module div_32_5(X, Q);//, R );

input  [32:1] X;
output [30:1] Q;  
//output [3:1] R;  


wire [8:1] r_1;
wire [8:1] r_2;
wire [8:1] r_3;
wire [7:1] r_4;
wire [6:1] r_5;

wire [5:1] sum_res;
wire [3:1] sum;

wire [10:1] q_1;
wire [16:1] q_2;
wire [22:1] q_3;
wire [28:1] q_4;
wire [33:1] q_5;


q_1 label1 ( .x0(X[9]),.x1(X[8]),.x2(X[7]),.x3(X[6]),.x4(X[5]),.x5(X[4]),
.z0(q_1[10]),.z1(q_1[9]),.z2(q_1[8]),.z3(q_1[7]),.z4(q_1[6]),.z5(q_1[5]),.z6(q_1[4]),.z7(q_1[3]),.z8(q_1[2]),.z9(q_1[1]));

q_2 label2 ( .x0(X[15]),.x1(X[14]),.x2(X[13]),.x3(X[12]),.x4(X[11]),.x5(X[10]),
.z00(q_2[16]),.z01(q_2[15]),.z02(q_2[14]),.z03(q_2[13]),.z04(q_2[12]),.z05(q_2[11]),.z06(q_2[10]),.z07(q_2[9]),.z08(q_2[8]),.z09(q_2[7]),.z10(q_2[6]),.z11(q_2[5]),.z12(q_2[4]),.z13(q_2[3]),.z14(q_2[2]),.z15(q_2[1]));

q_3 label3 ( .x0(X[21]),.x1(X[20]),.x2(X[19]),.x3(X[18]),.x4(X[17]),.x5(X[16]),
.z00(q_3[22]),.z01(q_3[21]),.z02(q_3[20]),.z03(q_3[19]),.z04(q_3[18]),.z05(q_3[17]),.z06(q_3[16]),.z07(q_3[15]),.z08(q_3[14]),.z09(q_3[13]),.z10(q_3[12]),.z11(q_3[11]),.z12(q_3[10]),.z13(q_3[9]),.z14(q_3[8]),.z15(q_3[7]),.z16(q_3[6]),.z17(q_3[5]),.z18(q_3[4]),.z19(q_3[3]),.z20(q_3[2]),.z21(q_3[1]));

q_4 label4 ( .x0(X[27]),.x1(X[26]),.x2(X[25]),.x3(X[24]),.x4(X[23]),.x5(X[22]),
.z00(q_4[28]),.z01(q_4[27]),.z02(q_4[26]),.z03(q_4[25]),.z04(q_4[24]),.z05(q_4[23]),.z06(q_4[22]),.z07(q_4[21]),.z08(q_4[20]),.z09(q_4[19]),.z10(q_4[18]),.z11(q_4[17]),.z12(q_4[16]),.z13(q_4[15]),.z14(q_4[14]),.z15(q_4[13]),.z16(q_4[12]),.z17(q_4[11]),.z18(q_4[10]),.z19(q_4[9]),.z20(q_4[8]),.z21(q_4[7]),.z22(q_4[6]),.z23(q_4[5]),.z24(q_4[4]),.z25(q_4[3]),.z26(q_4[2]),.z27(q_4[1]));

q_5 label5 ( .x0(X[32]),.x1(X[31]),.x2(X[30]),.x3(X[29]),.x4(X[28]),
.z00(q_5[33]),.z01(q_5[32]),.z02(q_5[31]),.z03(q_5[30]),.z04(q_5[29]),.z05(q_5[28]),.z06(q_5[27]),.z07(q_5[26]),.z08(q_5[25]),.z09(q_5[24]),.z10(q_5[23]),.z11(q_5[22]),.z12(q_5[21]),.z13(q_5[20]),.z14(q_5[19]),.z15(q_5[18]),.z16(q_5[17]),.z17(q_5[16]),.z18(q_5[15]),.z19(q_5[14]),.z20(q_5[13]),.z21(q_5[12]),.z22(q_5[11]),.z23(q_5[10]),.z24(q_5[9]),.z25(q_5[8]),.z26(q_5[7]),.z27(q_5[6]),.z28(q_5[5]),.z29(q_5[4]),.z30(q_5[3]),.z31(q_5[2]),.z32(q_5[1]));


assign sum_res = X[3:1] + q_1[3:1] + q_2[3:1] + q_3[3:1]+ q_4[3:1]+ q_5[3:1];

quot  label10 (.x0(sum_res[5]),.x1(sum_res[4]),.x2(sum_res[3]),.x3(sum_res[2]),.x4(sum_res[1]),
                  .z0(sum[3]),.z1(sum[2]),.z2(sum[1]));

assign r_1 = q_1[9:4] + q_2[9:4] + q_3[9:4]+ q_4[9:4] + q_5[9:4];

assign r_2 = r_1[8:7] + q_1[10] + q_2[15:10] + q_3[15:10] + q_4[15:10] + q_5[15:10];

assign r_3 = r_2[8:7] + q_2[16] + q_3[21:16] + q_4[21:16] + q_5[21:16];

assign r_4 = r_3[8:7] + q_3[22] + q_4[27:22] + q_5[27:22];

assign r_5 = r_4[7] + q_4[28] + q_5[33:28];


assign Q = {r_5[6:1], r_4[6:1], r_3[6:1], r_2[6:1], r_1[6:1]} + sum;


endmodule