module div_64_11(X, R);//, R );

input  [64:1] X;
//output [61:1] Q;  
output [4:1] R;  

wire [7:1] sum_res;

wire [4:1] q_1;
wire [4:1] q_2;
wire [4:1] q_3;
wire [4:1] q_4;
wire [4:1] q_5;
wire [4:1] q_6;
wire [4:1] q_7;
wire [4:1] q_8;
wire [4:1] q_9;
wire [4:1] q_10;


q_1 label1 ( .x0(X[10]),.x1(X[9]),.x2(X[8]),.x3(X[7]),.x4(X[6]),.x5(X[5]),
.z0(q_1[4]),.z1(q_1[3]),.z2(q_1[2]),.z3(q_1[1]));

q_2 label2 ( .x0(X[16]),.x1(X[15]),.x2(X[14]),.x3(X[13]),.x4(X[12]),.x5(X[11]),
.z0(q_2[4]),.z1(q_2[3]),.z2(q_2[2]),.z3(q_2[1]));

q_3 label3 ( .x0(X[22]),.x1(X[21]),.x2(X[20]),.x3(X[19]),.x4(X[18]),.x5(X[17]),
.z0(q_3[4]),.z1(q_3[3]),.z2(q_3[2]),.z3(q_3[1]));

q_4 label4 ( .x0(X[28]),.x1(X[27]),.x2(X[26]),.x3(X[25]),.x4(X[24]),.x5(X[23]),
.z0(q_4[4]),.z1(q_4[3]),.z2(q_4[2]),.z3(q_4[1]));

q_5 label5 ( .x0(X[34]),.x1(X[33]),.x2(X[32]),.x3(X[31]),.x4(X[30]),.x5(X[29]),
.z0(q_5[4]),.z1(q_5[3]),.z2(q_5[2]),.z3(q_5[1]));

q_6 label6 ( .x0(X[40]),.x1(X[39]),.x2(X[38]),.x3(X[37]),.x4(X[36]),.x5(X[35]),
.z0(q_6[4]),.z1(q_6[3]),.z2(q_6[2]),.z3(q_6[1]));

q_7 label7 ( .x0(X[46]),.x1(X[45]),.x2(X[44]),.x3(X[43]),.x4(X[42]),.x5(X[41]),
.z0(q_7[4]),.z1(q_7[3]),.z2(q_7[2]),.z3(q_7[1]));

q_8 label8 ( .x0(X[52]),.x1(X[51]),.x2(X[50]),.x3(X[49]),.x4(X[48]),.x5(X[47]),
.z0(q_8[4]),.z1(q_8[3]),.z2(q_8[2]),.z3(q_8[1]));

q_9 label9 ( .x0(X[58]),.x1(X[57]),.x2(X[56]),.x3(X[55]),.x4(X[54]),.x5(X[53]),
.z0(q_9[4]),.z1(q_9[3]),.z2(q_9[2]),.z3(q_9[1]));

q_10 label10 ( .x0(X[64]),.x1(X[63]),.x2(X[62]),.x3(X[61]),.x4(X[60]),.x5(X[59]),
.z0(q_10[4]),.z1(q_10[3]),.z2(q_10[2]),.z3(q_10[1]));

assign sum_res = X[4:1] + q_1[4:1] + q_2[4:1] + q_3[4:1] + q_4[4:1] + q_5[4:1] + q_6[4:1] + q_7[4:1] + q_8[4:1] + q_9[4:1] + q_10[4:1];

res  label12 (.x0(sum_res[7]),.x1(sum_res[6]),.x2(sum_res[5]),.x3(sum_res[4]),.x4(sum_res[3]),.x5(sum_res[2]),.x6(sum_res[1]),
          .z0(R[4]),.z1(R[3]),.z2(R[2]),.z3(R[1]));


endmodule