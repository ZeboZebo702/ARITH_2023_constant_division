module div_32_11(X, Q, R );

input  [32:1] X;
output [29:1] Q;  
output [4:1] R;  

wire [8:1] r_1;
wire [8:1] r_2;
wire [8:1] r_3;
wire [7:1] r_4;
wire [5:1] r_5;

wire [6:1] sum_res;
wire [7:1] sum;

wire [11:1] q_1;
wire [17:1] q_2;
wire [23:1] q_3;
wire [29:1] q_4;
wire [33:1] q_5;


q_1 label1 ( .x0(X[10]),.x1(X[9]),.x2(X[8]),.x3(X[7]),.x4(X[6]),.x5(X[5]),
.z00(q_1[11]),.z01(q_1[10]),.z02(q_1[9]),.z03(q_1[8]),.z04(q_1[7]),.z05(q_1[6]),.z06(q_1[5]),.z07(q_1[4]),.z08(q_1[3]),.z09(q_1[2]),.z10(q_1[1]));

q_2 label2 ( .x0(X[16]),.x1(X[15]),.x2(X[14]),.x3(X[13]),.x4(X[12]),.x5(X[11]),
.z00(q_2[17]),.z01(q_2[16]),.z02(q_2[15]),.z03(q_2[14]),.z04(q_2[13]),.z05(q_2[12]),.z06(q_2[11]),.z07(q_2[10]),.z08(q_2[9]),.z09(q_2[8]),.z10(q_2[7]),.z11(q_2[6]),.z12(q_2[5]),.z13(q_2[4]),.z14(q_2[3]),.z15(q_2[2]),.z16(q_2[1]));

q_3 label3 ( .x0(X[22]),.x1(X[21]),.x2(X[20]),.x3(X[19]),.x4(X[18]),.x5(X[17]),
.z00(q_3[23]),.z01(q_3[22]),.z02(q_3[21]),.z03(q_3[20]),.z04(q_3[19]),.z05(q_3[18]),.z06(q_3[17]),.z07(q_3[16]),.z08(q_3[15]),.z09(q_3[14]),.z10(q_3[13]),.z11(q_3[12]),.z12(q_3[11]),.z13(q_3[10]),.z14(q_3[9]),.z15(q_3[8]),.z16(q_3[7]),.z17(q_3[6]),.z18(q_3[5]),.z19(q_3[4]),.z20(q_3[3]),.z21(q_3[2]),.z22(q_3[1]));

q_4 label4 ( .x0(X[28]),.x1(X[27]),.x2(X[26]),.x3(X[25]),.x4(X[24]),.x5(X[23]),
.z00(q_4[29]),.z01(q_4[28]),.z02(q_4[27]),.z03(q_4[26]),.z04(q_4[25]),.z05(q_4[24]),.z06(q_4[23]),.z07(q_4[22]),.z08(q_4[21]),.z09(q_4[20]),.z10(q_4[19]),.z11(q_4[18]),.z12(q_4[17]),.z13(q_4[16]),.z14(q_4[15]),.z15(q_4[14]),.z16(q_4[13]),.z17(q_4[12]),.z18(q_4[11]),.z19(q_4[10]),.z20(q_4[9]),.z21(q_4[8]),.z22(q_4[7]),.z23(q_4[6]),.z24(q_4[5]),.z25(q_4[4]),.z26(q_4[3]),.z27(q_4[2]),.z28(q_4[1]));

q_5 label5 ( .x0(X[32]),.x1(X[31]),.x2(X[30]),.x3(X[29]),
.z00(q_5[33]),.z01(q_5[32]),.z02(q_5[31]),.z03(q_5[30]),.z04(q_5[29]),.z05(q_5[28]),.z06(q_5[27]),.z07(q_5[26]),.z08(q_5[25]),.z09(q_5[24]),.z10(q_5[23]),.z11(q_5[22]),.z12(q_5[21]),.z13(q_5[20]),.z14(q_5[19]),.z15(q_5[18]),.z16(q_5[17]),.z17(q_5[16]),.z18(q_5[15]),.z19(q_5[14]),.z20(q_5[13]),.z21(q_5[12]),.z22(q_5[11]),.z23(q_5[10]),.z24(q_5[9]),.z25(q_5[8]),.z26(q_5[7]),.z27(q_5[6]),.z28(q_5[5]),.z29(q_5[4]),.z30(q_5[3]),.z31(q_5[2]),.z32(q_5[1]));


assign sum_res = X[4:1] + q_1[4:1] + q_2[4:1] + q_3[4:1] + q_4[4:1] + q_5[4:1];

quot_res  label6 (.x0(sum_res[6]),.x1(sum_res[5]),.x2(sum_res[4]),.x3(sum_res[3]),.x4(sum_res[2]),.x5(sum_res[1]),
          .z0(sum[7]),.z1(sum[6]),.z2(sum[5]),.z3(sum[4]),.z4(sum[3]),.z5(sum[2]),.z6(sum[1]));

assign r_1 = q_1[10:5] + q_2[10:5] + q_3[10:5] + q_4[10:5] + q_5[10:5];

assign r_2 = r_1[8:7] + q_1[11] + q_2[16:11]+ q_3[16:11]+ q_4[16:11]+ q_5[16:11];

assign r_3 = r_2[8:7] + q_2[17] + q_3[22:17]+ q_4[22:17]+ q_5[22:17];

assign r_4 = r_3[8:7] + q_3[23]+ q_4[28:23]+ q_5[28:23];

assign r_5 = r_4[7] + q_4[29]+ q_5[33:29];



assign Q = {r_5, r_4[6:1], r_3[6:1], r_2[6:1], r_1[6:1]} + sum[7:5];

assign R = sum[4:1];

endmodule