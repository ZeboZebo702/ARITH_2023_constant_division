module div_32_23(X, Q, R );

input  [32:1] X;
output [28:1] Q;  
output [5:1] R;  

wire [28:1] Q_temp;

wire [9:1] r_1;
wire [8:1] r_2;
wire [8:1] r_3;
wire [7:1] r_4;
wire [4:1] r_5;

wire [7:1] sum_res;
wire [8:1] sum;

wire [12:1] q_1;
wire [18:1] q_2;
wire [24:1] q_3;
wire [30:1] q_4;
wire [33:1] q_5;

q_1 label1 ( .x0(X[11]),.x1(X[10]),.x2(X[9]),.x3(X[8]),.x4(X[7]),.x5(X[6]),
.z00(q_1[12]),.z01(q_1[11]),.z02(q_1[10]),.z03(q_1[9]),.z04(q_1[8]),.z05(q_1[7]),.z06(q_1[6]),.z07(q_1[5]),.z08(q_1[4]),.z09(q_1[3]),.z10(q_1[2]),.z11(q_1[1]));

q_2 label2 ( .x0(X[17]),.x1(X[16]),.x2(X[15]),.x3(X[14]),.x4(X[13]),.x5(X[12]),
.z00(q_2[18]),.z01(q_2[17]),.z02(q_2[16]),.z03(q_2[15]),.z04(q_2[14]),.z05(q_2[13]),.z06(q_2[12]),.z07(q_2[11]),.z08(q_2[10]),.z09(q_2[9]),.z10(q_2[8]),.z11(q_2[7]),.z12(q_2[6]),.z13(q_2[5]),.z14(q_2[4]),.z15(q_2[3]),.z16(q_2[2]),.z17(q_2[1]));

q_3 label3 ( .x0(X[23]),.x1(X[22]),.x2(X[21]),.x3(X[20]),.x4(X[19]),.x5(X[18]),
.z00(q_3[24]),.z01(q_3[23]),.z02(q_3[22]),.z03(q_3[21]),.z04(q_3[20]),.z05(q_3[19]),.z06(q_3[18]),.z07(q_3[17]),.z08(q_3[16]),.z09(q_3[15]),.z10(q_3[14]),.z11(q_3[13]),.z12(q_3[12]),.z13(q_3[11]),.z14(q_3[10]),.z15(q_3[9]),.z16(q_3[8]),.z17(q_3[7]),.z18(q_3[6]),.z19(q_3[5]),.z20(q_3[4]),.z21(q_3[3]),.z22(q_3[2]),.z23(q_3[1]));

q_4 label4 ( .x0(X[29]),.x1(X[28]),.x2(X[27]),.x3(X[26]),.x4(X[25]),.x5(X[24]),
.z00(q_4[30]),.z01(q_4[29]),.z02(q_4[28]),.z03(q_4[27]),.z04(q_4[26]),.z05(q_4[25]),.z06(q_4[24]),.z07(q_4[23]),.z08(q_4[22]),.z09(q_4[21]),.z10(q_4[20]),.z11(q_4[19]),.z12(q_4[18]),.z13(q_4[17]),.z14(q_4[16]),.z15(q_4[15]),.z16(q_4[14]),.z17(q_4[13]),.z18(q_4[12]),.z19(q_4[11]),.z20(q_4[10]),.z21(q_4[9]),.z22(q_4[8]),.z23(q_4[7]),.z24(q_4[6]),.z25(q_4[5]),.z26(q_4[4]),.z27(q_4[3]),.z28(q_4[2]),.z29(q_4[1]));

q_5 label5 ( .x0(X[32]),.x1(X[31]),.x2(X[30]),
.z00(q_5[33]),.z01(q_5[32]),.z02(q_5[31]),.z03(q_5[30]),.z04(q_5[29]),.z05(q_5[28]),.z06(q_5[27]),.z07(q_5[26]),.z08(q_5[25]),.z09(q_5[24]),.z10(q_5[23]),.z11(q_5[22]),.z12(q_5[21]),.z13(q_5[20]),.z14(q_5[19]),.z15(q_5[18]),.z16(q_5[17]),.z17(q_5[16]),.z18(q_5[15]),.z19(q_5[14]),.z20(q_5[13]),.z21(q_5[12]),.z22(q_5[11]),.z23(q_5[10]),.z24(q_5[9]),.z25(q_5[8]),.z26(q_5[7]),.z27(q_5[6]),.z28(q_5[5]),.z29(q_5[4]),.z30(q_5[3]),.z31(q_5[2]),.z32(q_5[1]));


assign sum_res = X[5:1] + q_1[5:1] + q_2[5:1] + q_3[5:1] + q_4[5:1] + q_5[5:1];

quot_res  label10 (.x0(sum_res[7]),.x1(sum_res[6]),.x2(sum_res[5]),.x3(sum_res[4]),.x4(sum_res[3]),
		  .x5(sum_res[2]),.x6(sum_res[1]),
                  .z0(sum[8]),.z1(sum[7]),.z2(sum[6]),.z3(sum[5]),.z4(sum[4]),
		  .z5(sum[3]),.z6(sum[2]),.z7(sum[1]));


assign r_1 = q_1[11:6] + q_2[11:6] + q_3[11:6] + q_4[11:6] + q_5[11:6];

assign r_2 = r_1[9:7] + q_1[12] + q_2[17:12] + q_3[17:12] + q_4[17:12] + q_5[17:12];

assign r_3 = r_2[8:7] + q_2[18] + q_3[23:18] + q_4[23:18] + q_5[23:18];

assign r_4 = r_3[8:7] + q_3[24] + q_4[29:24] + q_5[29:24];

assign r_5 = r_4[7] + q_4[30] + q_5[33:30];

assign Q_temp = {r_5[4:1], r_4[6:1], r_3[6:1], r_2[6:1], r_1[6:1]};


assign Q = Q_temp + sum[8:6];

assign R = sum[5:1]; 

endmodule