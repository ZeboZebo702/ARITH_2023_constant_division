module div_64_5(X, R);//, R );

input  [64:1] X;
//output [62:1] Q;  
output [3:1] R;  



wire [6:1] sum_res;

wire [3:1] q_1;
wire [3:1] q_2;
wire [3:1] q_3;
wire [3:1] q_4;
wire [3:1] q_5;
wire [3:1] q_6;
wire [3:1] q_7;
wire [3:1] q_8;
wire [3:1] q_9;
wire [3:1] q_10;
wire [3:1] q_11;


q_1 label1 ( .x0(X[9]),.x1(X[8]),.x2(X[7]),.x3(X[6]),.x4(X[5]),.x5(X[4]),
.z0(q_1[3]),.z1(q_1[2]),.z2(q_1[1]));

q_2 label2 ( .x0(X[15]),.x1(X[14]),.x2(X[13]),.x3(X[12]),.x4(X[11]),.x5(X[10]),
.z0(q_2[3]),.z1(q_2[2]),.z2(q_2[1]));

q_3 label3 ( .x0(X[21]),.x1(X[20]),.x2(X[19]),.x3(X[18]),.x4(X[17]),.x5(X[16]),
.z0(q_3[3]),.z1(q_3[2]),.z2(q_3[1]));

q_4 label4 ( .x0(X[27]),.x1(X[26]),.x2(X[25]),.x3(X[24]),.x4(X[23]),.x5(X[22]),
.z0(q_4[3]),.z1(q_4[2]),.z2(q_4[1]));

q_5 label5 ( .x0(X[33]),.x1(X[32]),.x2(X[31]),.x3(X[30]),.x4(X[29]),.x5(X[28]),
.z0(q_5[3]),.z1(q_5[2]),.z2(q_5[1]));

q_6 label6 ( .x0(X[39]),.x1(X[38]),.x2(X[37]),.x3(X[36]),.x4(X[35]),.x5(X[34]),
.z0(q_6[3]),.z1(q_6[2]),.z2(q_6[1]));

q_7 label7 ( .x0(X[45]),.x1(X[44]),.x2(X[43]),.x3(X[42]),.x4(X[41]),.x5(X[40]),
.z0(q_7[3]),.z1(q_7[2]),.z2(q_7[1]));

q_8 label8 ( .x0(X[51]),.x1(X[50]),.x2(X[49]),.x3(X[48]),.x4(X[47]),.x5(X[46]),
.z0(q_8[3]),.z1(q_8[2]),.z2(q_8[1]));

q_9 label9 ( .x0(X[57]),.x1(X[56]),.x2(X[55]),.x3(X[54]),.x4(X[53]),.x5(X[52]),
.z0(q_9[3]),.z1(q_9[2]),.z2(q_9[1]));

q_10 label10 ( .x0(X[63]),.x1(X[62]),.x2(X[61]),.x3(X[60]),.x4(X[59]),.x5(X[58]),
.z0(q_10[3]),.z1(q_10[2]),.z2(q_10[1]));

q_11 label11 ( .x0(X[64]),
.z0(q_11[3]),.z1(q_11[2]),.z2(q_11[1]));


assign sum_res = X[3:1] + q_1[3:1] + q_2[3:1] + q_3[3:1]+ q_4[3:1]+ q_5[3:1] + q_6[3:1] + q_7[3:1] + q_8[3:1]+ q_9[3:1]+ q_10[3:1] + q_11[3:1];

res  label12 (.x0(sum_res[6]),.x1(sum_res[5]),.x2(sum_res[4]),.x3(sum_res[3]),.x4(sum_res[2]),.x5(sum_res[1]),
                  .z0(R[3]),.z1(R[2]),.z2(R[1]));


endmodule