module div_64_23(X, R );

input  [64:1] X;
//output [28:1] Q;  
output [5:1] R;  

//wire [28:1] Q_temp;

wire [5:1] r_1;
wire [5:1] r_2;
wire [5:1] r_3;
wire [5:1] r_4;
wire [5:1] r_5;
wire [5:1] q_6;
wire [5:1] q_7;
wire [5:1] q_8;
wire [5:1] q_9;
wire [5:1] q_10;

//wire [7:1] sum_res;
wire [8:1] res;


q_1 label1 (.x0(X[11]),.x1(X[10]),.x2(X[9]),.x3(X[8]),.x4(X[7]),.x5(X[6]),
.z0(r_1[5]),.z1(r_1[4]),.z2(r_1[3]),.z3(r_1[2]),.z4(r_1[1]));

q_2 label2 ( .x0(X[17]),.x1(X[16]),.x2(X[15]),.x3(X[14]),.x4(X[13]),.x5(X[12]),
.z0(r_2[5]),.z1(r_2[4]),.z2(r_2[3]),.z3(r_2[2]),.z4(r_2[1]));

q_3 label3 ( .x0(X[23]),.x1(X[22]),.x2(X[21]),.x3(X[20]),.x4(X[19]),.x5(X[18]),
.z0(r_3[5]),.z1(r_3[4]),.z2(r_3[3]),.z3(r_3[2]),.z4(r_3[1]));

q_4 label4 ( .x0(X[29]),.x1(X[28]),.x2(X[27]),.x3(X[26]),.x4(X[25]),.x5(X[24]),
.z0(r_4[5]),.z1(r_4[4]),.z2(r_4[3]),.z3(r_4[2]),.z4(r_4[1]));

q_5 label5 ( .x0(X[35]),.x1(X[34]),.x2(X[33]),.x3(X[32]),.x4(X[31]),.x5(X[30]),
.z0(r_5[5]),.z1(r_5[4]),.z2(r_5[3]),.z3(r_5[2]),.z4(r_5[1]));

q_6 label6 ( .x0(X[41]),.x1(X[40]),.x2(X[39]),.x3(X[38]),.x4(X[37]),.x5(X[36]),
.z0(q_6[5]),.z1(q_6[4]),.z2(q_6[3]),.z3(q_6[2]),.z4(q_6[1]));

q_7 label7 ( .x0(X[47]),.x1(X[46]),.x2(X[45]),.x3(X[44]),.x4(X[43]),.x5(X[42]),
.z0(q_7[5]),.z1(q_7[4]),.z2(q_7[3]),.z3(q_7[2]),.z4(q_7[1]));

q_8 label8 ( .x0(X[53]),.x1(X[52]),.x2(X[51]),.x3(X[50]),.x4(X[49]),.x5(X[48]),
.z0(q_8[5]),.z1(q_8[4]),.z2(q_8[3]),.z3(q_8[2]),.z4(q_8[1]));

q_9 label9 ( .x0(X[59]),.x1(X[58]),.x2(X[57]),.x3(X[56]),.x4(X[55]),.x5(X[54]),
.z0(q_9[5]),.z1(q_9[4]),.z2(q_9[3]),.z3(q_9[2]),.z4(q_9[1]));

q_10 label10 ( .x0(X[64]),.x1(X[63]),.x2(X[62]),.x3(X[61]),.x4(X[60]),
.z0(q_10[5]),.z1(q_10[4]),.z2(q_10[3]),.z3(q_10[2]),.z4(q_10[1])); 

assign res = X[5:1] + r_1 + r_2 + r_3 + r_4 + r_5 + q_6 + q_7 + q_8 + q_9 + q_10;

res  label11 (.x0(res[8]),.x1(res[7]),.x2(res[6]),.x3(res[5]),.x4(res[4]),.x5(res[3]),.x6(res[2]),.x7(res[1]),
                  .z0(R[5]),.z1(R[4]),.z2(R[3]),.z3(R[2]),.z4(R[1]));


endmodule