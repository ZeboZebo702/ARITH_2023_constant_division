module div_32_23(X, R );

input  [32:1] X;
//output [28:1] Q;  
output [5:1] R;  

//wire [28:1] Q_temp;

wire [5:1] r_1;
wire [5:1] r_2;
wire [5:1] r_3;
wire [5:1] r_4;
wire [5:1] r_5;

wire [7:1] sum_res;
//wire [8:1] res;


q_1 label1 (.x0(X[11]),.x1(X[10]),.x2(X[9]),.x3(X[8]),.x4(X[7]),.x5(X[6]),
.z0(r_1[5]),.z1(r_1[4]),.z2(r_1[3]),.z3(r_1[2]),.z4(r_1[1]));

q_2 label2 ( .x0(X[17]),.x1(X[16]),.x2(X[15]),.x3(X[14]),.x4(X[13]),.x5(X[12]),
.z0(r_2[5]),.z1(r_2[4]),.z2(r_2[3]),.z3(r_2[2]),.z4(r_2[1]));

q_3 label3 ( .x0(X[23]),.x1(X[22]),.x2(X[21]),.x3(X[20]),.x4(X[19]),.x5(X[18]),
.z0(r_3[5]),.z1(r_3[4]),.z2(r_3[3]),.z3(r_3[2]),.z4(r_3[1]));

q_4 label4 ( .x0(X[29]),.x1(X[28]),.x2(X[27]),.x3(X[26]),.x4(X[25]),.x5(X[24]),
.z0(r_4[5]),.z1(r_4[4]),.z2(r_4[3]),.z3(r_4[2]),.z4(r_4[1]));

q_5 label5 ( .x0(X[32]),.x1(X[31]),.x2(X[30]),
.z0(r_5[5]),.z1(r_5[4]),.z2(r_5[3]),.z3(r_5[2]),.z4(r_5[1]));


assign sum_res = X[5:1] + r_1 + r_2 + r_3 + r_4 + r_5;

res  label10 (.x0(sum_res[7]),.x1(sum_res[6]),.x2(sum_res[5]),.x3(sum_res[4]),.x4(sum_res[3]),
		  .x5(sum_res[2]),.x6(sum_res[1]),
                  .z0(R[5]),.z1(R[4]),.z2(R[3]),.z3(R[2]),.z4(R[1]));


endmodule