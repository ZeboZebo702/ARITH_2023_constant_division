// Benchmark "q_5" written by ABC on Mon Feb 27 04:09:45 2023

module q_5 ( 
    x0,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35  );
  input  x0;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35;
  assign z01 = 1'b0;
  assign z00 = x0;
  assign z02 = 1'b0;
  assign z03 = x0;
  assign z04 = 1'b0;
  assign z05 = 1'b0;
  assign z06 = 1'b0;
  assign z07 = 1'b0;
  assign z08 = x0;
  assign z09 = x0;
  assign z10 = x0;
  assign z11 = x0;
  assign z12 = x0;
  assign z13 = x0;
  assign z14 = 1'b0;
  assign z15 = x0;
  assign z16 = x0;
  assign z17 = 1'b0;
  assign z18 = x0;
  assign z19 = x0;
  assign z20 = x0;
  assign z21 = x0;
  assign z22 = 1'b0;
  assign z23 = 1'b0;
  assign z24 = 1'b0;
  assign z25 = 1'b0;
  assign z26 = 1'b0;
  assign z27 = 1'b0;
  assign z28 = x0;
  assign z29 = 1'b0;
  assign z30 = 1'b0;
  assign z31 = 1'b0;
  assign z32 = x0;
  assign z33 = x0;
  assign z34 = x0;
  assign z35 = x0;
endmodule


