module div_24_47(X, Q, R );

input  [24:1] X;
output [19:1] Q;  
output [6:1] R;  

wire [19:1] Q_tmp;
wire [8:1] r_1;
wire [7:1] r_2;
wire [6:1] r_3;
wire r_4;

wire [8:1] sum_res;
wire [8:1] sum;

wire [13:1] q_1;
wire [19:1] q_2;
wire [25:1] q_3;

q_1  label1 (.x0(X[12]),.x1(X[11]),.x2(X[10]),.x3(X[9]),.x4(X[8]),.x5(X[7]),
          .z00(q_1[13]),.z01(q_1[12]),.z02(q_1[11]),.z03(q_1[10]),.z04(q_1[9]),.z05(q_1[8]),.z06(q_1[7]),.z07(q_1[6]),
	  .z08(q_1[5]),.z09(q_1[4]),.z10(q_1[3]),.z11(q_1[2]),.z12(q_1[1]));

q_2  label2 (.x0(X[18]),.x1(X[17]),.x2(X[16]),.x3(X[15]),.x4(X[14]),.x5(X[13]),
	  .z00(q_2[19]),.z01(q_2[18]),.z02(q_2[17]),.z03(q_2[16]),.z04(q_2[15]),	
      .z05(q_2[14]),.z06(q_2[13]),.z07(q_2[12]),.z08(q_2[11]),.z09(q_2[10]),.z10(q_2[9]),
	  .z11(q_2[8]),.z12(q_2[7]),.z13(q_2[6]),.z14(q_2[5]),.z15(q_2[4]),.z16(q_2[3]),.z17(q_2[2]),.z18(q_2[1]));

q_3  label3 (.x0(X[24]),.x1(X[23]),.x2(X[22]),.x3(X[21]),.x4(X[20]),.x5(X[19]),
	  .z00(q_3[25]),.z01(q_3[24]),.z02(q_3[23]),.z03(q_3[22]),.z04(q_3[21]),
      .z05(q_3[20]),.z06(q_3[19]),.z07(q_3[18]),.z08(q_3[17]),.z09(q_3[16]),.z10(q_3[15]),
	  .z11(q_3[14]),.z12(q_3[13]),.z13(q_3[12]),.z14(q_3[11]),.z15(q_3[10]),
	  .z16(q_3[9]),.z17(q_3[8]),.z18(q_3[7]),.z19(q_3[6]),.z20(q_3[5]),.z21(q_3[4]),.z22(q_3[3]),.z23(q_3[2]),.z24(q_3[1]));

assign sum_res = X[6:1] + q_1[6:1] + q_2[6:1] + q_3[6:1];

quot_res  label4 (.x0(sum_res[8]),.x1(sum_res[7]),.x2(sum_res[6]),.x3(sum_res[5]),.x4(sum_res[4]),.x5(sum_res[3]),.x6(sum_res[2]),.x7(sum_res[1]),
          .z0(sum[8]),.z1(sum[7]),.z2(sum[6]),.z3(sum[5]),.z4(sum[4]),.z5(sum[3]),.z6(sum[2]),.z7(sum[1]));

assign r_1 = q_1[12:7] + q_2[12:7] + q_3[12:7];

assign r_2 = r_1[8:7] + q_1[13] + q_2[18:13] + q_3[18:13];

assign r_3 = r_2[7] + q_2[19] + q_3[24:19];

assign r_4 = q_3[25];

assign Q_tmp = {r_4, r_3[6:1], r_2[6:1], r_1[6:1]};

assign Q = Q_tmp + sum[8:7];

assign R = sum[6:1];

endmodule