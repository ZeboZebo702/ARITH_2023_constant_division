// Benchmark "q_11" written by ABC on Tue Jul 11 01:01:40 2023

module q_11 ( 
    x0,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63  );
  input  x0;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63;
  assign z00 = x0;
  assign z01 = x0;
  assign z02 = 1'b0;
  assign z03 = 1'b0;
  assign z04 = x0;
  assign z05 = x0;
  assign z06 = 1'b0;
  assign z07 = 1'b0;
  assign z08 = x0;
  assign z09 = x0;
  assign z10 = 1'b0;
  assign z11 = 1'b0;
  assign z12 = x0;
  assign z13 = x0;
  assign z14 = 1'b0;
  assign z15 = 1'b0;
  assign z16 = x0;
  assign z17 = x0;
  assign z18 = 1'b0;
  assign z19 = 1'b0;
  assign z20 = x0;
  assign z21 = x0;
  assign z22 = 1'b0;
  assign z23 = 1'b0;
  assign z24 = x0;
  assign z25 = x0;
  assign z26 = 1'b0;
  assign z27 = 1'b0;
  assign z28 = x0;
  assign z29 = x0;
  assign z30 = 1'b0;
  assign z31 = 1'b0;
  assign z32 = x0;
  assign z33 = x0;
  assign z34 = 1'b0;
  assign z35 = 1'b0;
  assign z36 = x0;
  assign z37 = x0;
  assign z38 = 1'b0;
  assign z39 = 1'b0;
  assign z40 = x0;
  assign z41 = x0;
  assign z42 = 1'b0;
  assign z43 = 1'b0;
  assign z44 = x0;
  assign z45 = x0;
  assign z46 = 1'b0;
  assign z47 = 1'b0;
  assign z48 = x0;
  assign z49 = x0;
  assign z50 = 1'b0;
  assign z51 = 1'b0;
  assign z52 = x0;
  assign z53 = x0;
  assign z54 = 1'b0;
  assign z55 = 1'b0;
  assign z56 = x0;
  assign z57 = x0;
  assign z58 = 1'b0;
  assign z59 = 1'b0;
  assign z60 = x0;
  assign z61 = 1'b0;
  assign z62 = x0;
  assign z63 = x0;
endmodule


