module div_64_3(X, Q, R );

input  [64:1] X;
output [63:1] Q;  
output [2:1] R;  

wire [9:1] r_1;
wire [9:1] r_2;
wire [9:1] r_3;
wire [9:1] r_4;
wire [9:1] r_5;
wire [8:1] r_6;
wire [8:1] r_7;
wire [8:1] r_8;
wire [8:1] r_9;
wire [7:1] r_10;
wire [3:1] r_11;

wire [5:1] sum_res;
wire [6:1] sum;

wire [7:1] q_1;
wire [13:1] q_2;
wire [19:1] q_3;
wire [25:1] q_4;
wire [31:1] q_5;
wire [37:1] q_6;
wire [43:1] q_7;
wire [49:1] q_8;
wire [55:1] q_9;
wire [61:1] q_10;
wire [63:1] q_11;

q_1 label1 ( .x0(X[8]),.x1(X[7]),.x2(X[6]),.x3(X[5]),.x4(X[4]),.x5(X[3]),
.z0(q_1[7]),.z1(q_1[6]),.z2(q_1[5]),.z3(q_1[4]),.z4(q_1[3]),.z5(q_1[2]),.z6(q_1[1]));

q_2 label2 ( .x0(X[14]),.x1(X[13]),.x2(X[12]),.x3(X[11]),.x4(X[10]),.x5(X[9]),
.z00(q_2[13]),.z01(q_2[12]),.z02(q_2[11]),.z03(q_2[10]),.z04(q_2[9]),.z05(q_2[8]),.z06(q_2[7]),.z07(q_2[6]),.z08(q_2[5]),.z09(q_2[4]),.z10(q_2[3]),.z11(q_2[2]),.z12(q_2[1]));

q_3 label3 ( .x0(X[20]),.x1(X[19]),.x2(X[18]),.x3(X[17]),.x4(X[16]),.x5(X[15]),
.z00(q_3[19]),.z01(q_3[18]),.z02(q_3[17]),.z03(q_3[16]),.z04(q_3[15]),.z05(q_3[14]),.z06(q_3[13]),.z07(q_3[12]),.z08(q_3[11]),.z09(q_3[10]),.z10(q_3[9]),.z11(q_3[8]),.z12(q_3[7]),.z13(q_3[6]),.z14(q_3[5]),.z15(q_3[4]),.z16(q_3[3]),.z17(q_3[2]),.z18(q_3[1]));

q_4 label4 ( .x0(X[26]),.x1(X[25]),.x2(X[24]),.x3(X[23]),.x4(X[22]),.x5(X[21]),
.z00(q_4[25]),.z01(q_4[24]),.z02(q_4[23]),.z03(q_4[22]),.z04(q_4[21]),.z05(q_4[20]),.z06(q_4[19]),.z07(q_4[18]),.z08(q_4[17]),.z09(q_4[16]),.z10(q_4[15]),.z11(q_4[14]),.z12(q_4[13]),.z13(q_4[12]),.z14(q_4[11]),.z15(q_4[10]),.z16(q_4[9]),.z17(q_4[8]),.z18(q_4[7]),.z19(q_4[6]),.z20(q_4[5]),.z21(q_4[4]),.z22(q_4[3]),.z23(q_4[2]),.z24(q_4[1]));

q_5 label5 ( .x0(X[32]),.x1(X[31]),.x2(X[30]),.x3(X[29]),.x4(X[28]),.x5(X[27]),
.z00(q_5[31]),.z01(q_5[30]),.z02(q_5[29]),.z03(q_5[28]),.z04(q_5[27]),.z05(q_5[26]),.z06(q_5[25]),.z07(q_5[24]),.z08(q_5[23]),.z09(q_5[22]),.z10(q_5[21]),.z11(q_5[20]),.z12(q_5[19]),.z13(q_5[18]),.z14(q_5[17]),.z15(q_5[16]),.z16(q_5[15]),.z17(q_5[14]),.z18(q_5[13]),.z19(q_5[12]),.z20(q_5[11]),.z21(q_5[10]),.z22(q_5[9]),.z23(q_5[8]),.z24(q_5[7]),.z25(q_5[6]),.z26(q_5[5]),.z27(q_5[4]),.z28(q_5[3]),.z29(q_5[2]),.z30(q_5[1]));


q_6 label6 ( .x0(X[38]),.x1(X[37]),.x2(X[36]),.x3(X[35]),.x4(X[34]),.x5(X[33]),
.z00(q_6[37]),.z01(q_6[36]),.z02(q_6[35]),.z03(q_6[34]),.z04(q_6[33]),.z05(q_6[32]),.z06(q_6[31]),.z07(q_6[30]),.z08(q_6[29]),.z09(q_6[28]),
.z10(q_6[27]),.z11(q_6[26]),.z12(q_6[25]),.z13(q_6[24]),.z14(q_6[23]),.z15(q_6[22]),.z16(q_6[21]),.z17(q_6[20]),.z18(q_6[19]),.z19(q_6[18]),
.z20(q_6[17]),.z21(q_6[16]),.z22(q_6[15]),.z23(q_6[14]),.z24(q_6[13]),.z25(q_6[12]),.z26(q_6[11]),.z27(q_6[10]),.z28(q_6[9]),.z29(q_6[8]),
.z30(q_6[7]),.z31(q_6[6]),.z32(q_6[5]),.z33(q_6[4]),.z34(q_6[3]),.z35(q_6[2]),.z36(q_6[1]));

q_7 label7 ( .x0(X[44]),.x1(X[43]),.x2(X[42]),.x3(X[41]),.x4(X[40]),.x5(X[39]),
.z00(q_7[43]),.z01(q_7[42]),.z02(q_7[41]),.z03(q_7[40]),.z04(q_7[39]),.z05(q_7[38]),.z06(q_7[37]),.z07(q_7[36]),.z08(q_7[35]),.z09(q_7[34]),
.z10(q_7[33]),.z11(q_7[32]),.z12(q_7[31]),.z13(q_7[30]),.z14(q_7[29]),.z15(q_7[28]),.z16(q_7[27]),.z17(q_7[26]),.z18(q_7[25]),.z19(q_7[24]),
.z20(q_7[23]),.z21(q_7[22]),.z22(q_7[21]),.z23(q_7[20]),.z24(q_7[19]),.z25(q_7[18]),.z26(q_7[17]),.z27(q_7[16]),.z28(q_7[15]),.z29(q_7[14]),
.z30(q_7[13]),.z31(q_7[12]),.z32(q_7[11]),.z33(q_7[10]),.z34(q_7[9]),.z35(q_7[8]),.z36(q_7[7]),.z37(q_7[6]),.z38(q_7[5]),.z39(q_7[4]),
.z40(q_7[3]),.z41(q_7[2]),.z42(q_7[1]));

q_8 label8 ( .x0(X[50]),.x1(X[49]),.x2(X[48]),.x3(X[47]),.x4(X[46]),.x5(X[45]),
.z00(q_8[49]),.z01(q_8[48]),.z02(q_8[47]),.z03(q_8[46]),.z04(q_8[45]),.z05(q_8[44]),.z06(q_8[43]),.z07(q_8[42]),.z08(q_8[41]),.z09(q_8[40]),
.z10(q_8[39]),.z11(q_8[38]),.z12(q_8[37]),.z13(q_8[36]),.z14(q_8[35]),.z15(q_8[34]),.z16(q_8[33]),.z17(q_8[32]),.z18(q_8[31]),.z19(q_8[30]),
.z20(q_8[29]),.z21(q_8[28]),.z22(q_8[27]),.z23(q_8[26]),.z24(q_8[25]),.z25(q_8[24]),.z26(q_8[23]),.z27(q_8[22]),.z28(q_8[21]),.z29(q_8[20]),
.z30(q_8[19]),.z31(q_8[18]),.z32(q_8[17]),.z33(q_8[16]),.z34(q_8[15]),.z35(q_8[14]),.z36(q_8[13]),.z37(q_8[12]),.z38(q_8[11]),.z39(q_8[10]),
.z40(q_8[9]),.z41(q_8[8]),.z42(q_8[7]),.z43(q_8[6]),.z44(q_8[5]),.z45(q_8[4]),.z46(q_8[3]),.z47(q_8[2]),.z48(q_8[1]));

q_9 label9 ( .x0(X[56]),.x1(X[55]),.x2(X[54]),.x3(X[53]),.x4(X[52]),.x5(X[51]),
.z00(q_9[55]),.z01(q_9[54]),.z02(q_9[53]),.z03(q_9[52]),.z04(q_9[51]),.z05(q_9[50]),.z06(q_9[49]),.z07(q_9[48]),.z08(q_9[47]),.z09(q_9[46]),
.z10(q_9[45]),.z11(q_9[44]),.z12(q_9[43]),.z13(q_9[42]),.z14(q_9[41]),.z15(q_9[40]),.z16(q_9[39]),.z17(q_9[38]),.z18(q_9[37]),.z19(q_9[36]),
.z20(q_9[35]),.z21(q_9[34]),.z22(q_9[33]),.z23(q_9[32]),.z24(q_9[31]),.z25(q_9[30]),.z26(q_9[29]),.z27(q_9[28]),.z28(q_9[27]),.z29(q_9[26]),
.z30(q_9[25]),.z31(q_9[24]),.z32(q_9[23]),.z33(q_9[22]),.z34(q_9[21]),.z35(q_9[20]),.z36(q_9[19]),.z37(q_9[18]),.z38(q_9[17]),.z39(q_9[16]),
.z40(q_9[15]),.z41(q_9[14]),.z42(q_9[13]),.z43(q_9[12]),.z44(q_9[11]),.z45(q_9[10]),.z46(q_9[9]),.z47(q_9[8]),.z48(q_9[7]),.z49(q_9[6]),
.z50(q_9[5]),.z51(q_9[4]),.z52(q_9[3]),.z53(q_9[2]),.z54(q_9[1]));

q_10 label10 ( .x0(X[62]),.x1(X[61]),.x2(X[60]),.x3(X[59]),.x4(X[58]),.x5(X[57]),
.z00(q_10[61]),.z01(q_10[60]),.z02(q_10[59]),.z03(q_10[58]),.z04(q_10[57]),.z05(q_10[56]),.z06(q_10[55]),.z07(q_10[54]),.z08(q_10[53]),.z09(q_10[52]),
.z10(q_10[51]),.z11(q_10[50]),.z12(q_10[49]),.z13(q_10[48]),.z14(q_10[47]),.z15(q_10[46]),.z16(q_10[45]),.z17(q_10[44]),.z18(q_10[43]),.z19(q_10[42]),
.z20(q_10[41]),.z21(q_10[40]),.z22(q_10[39]),.z23(q_10[38]),.z24(q_10[37]),.z25(q_10[36]),.z26(q_10[35]),.z27(q_10[34]),.z28(q_10[33]),.z29(q_10[32]),
.z30(q_10[31]),.z31(q_10[30]),.z32(q_10[29]),.z33(q_10[28]),.z34(q_10[27]),.z35(q_10[26]),.z36(q_10[25]),.z37(q_10[24]),.z38(q_10[23]),.z39(q_10[22]),
.z40(q_10[21]),.z41(q_10[20]),.z42(q_10[19]),.z43(q_10[18]),.z44(q_10[17]),.z45(q_10[16]),.z46(q_10[15]),.z47(q_10[14]),.z48(q_10[13]),.z49(q_10[12]),
.z50(q_10[11]),.z51(q_10[10]),.z52(q_10[9]),.z53(q_10[8]),.z54(q_10[7]),.z55(q_10[6]),.z56(q_10[5]),.z57(q_10[4]),.z58(q_10[3]),.z59(q_10[2]),
.z60(q_10[1]));

q_11 label11 ( .x0(X[64]),.x1(X[63]),
.z00(q_11[63]),.z01(q_11[62]),.z02(q_11[61]),.z03(q_11[60]),.z04(q_11[59]),.z05(q_11[58]),.z06(q_11[57]),.z07(q_11[56]),.z08(q_11[55]),.z09(q_11[54]),
.z10(q_11[53]),.z11(q_11[52]),.z12(q_11[51]),.z13(q_11[50]),.z14(q_11[49]),.z15(q_11[48]),.z16(q_11[47]),.z17(q_11[46]),.z18(q_11[45]),.z19(q_11[44]),
.z20(q_11[43]),.z21(q_11[42]),.z22(q_11[41]),.z23(q_11[40]),.z24(q_11[39]),.z25(q_11[38]),.z26(q_11[37]),.z27(q_11[36]),.z28(q_11[35]),.z29(q_11[34]),
.z30(q_11[33]),.z31(q_11[32]),.z32(q_11[31]),.z33(q_11[30]),.z34(q_11[29]),.z35(q_11[28]),.z36(q_11[27]),.z37(q_11[26]),.z38(q_11[25]),.z39(q_11[24]),
.z40(q_11[23]),.z41(q_11[22]),.z42(q_11[21]),.z43(q_11[20]),.z44(q_11[19]),.z45(q_11[18]),.z46(q_11[17]),.z47(q_11[16]),.z48(q_11[15]),.z49(q_11[14]),
.z50(q_11[13]),.z51(q_11[12]),.z52(q_11[11]),.z53(q_11[10]),.z54(q_11[9]),.z55(q_11[8]),.z56(q_11[7]),.z57(q_11[6]),.z58(q_11[5]),.z59(q_11[4]),
.z60(q_11[3]),.z61(q_11[2]),.z62(q_11[1]));


assign sum_res = X[2:1] + q_1[2:1] + q_2[2:1] + q_3[2:1] + q_4[2:1] + q_5[2:1] +
		+ q_6[2:1] + q_7[2:1] + q_8[2:1] + q_9[2:1] + q_10[2:1] + q_11[2:1];

quot_res  label12 (.x0(sum_res[5]),.x1(sum_res[4]),.x2(sum_res[3]),.x3(sum_res[2]),.x4(sum_res[1]),
                  .z0(sum[6]),.z1(sum[5]),.z2(sum[4]),.z3(sum[3]),.z4(sum[2]),.z5(sum[1]));


assign r_1 = q_1[6:1] + q_2[6:1] + q_3[6:1] + q_4[6:1] + q_5[6:1] + q_6[6:1] + q_7[6:1] + q_8[6:1] + q_9[6:1] + q_10[6:1] + q_11[6:1];

assign r_2 = r_1[9:7] + q_1[7] + q_2[12:7] + q_3[12:7] + q_4[12:7] + q_5[12:7] + q_6[12:7] + q_7[12:7] + q_8[12:7] + q_9[12:7] + q_10[12:7] + q_11[12:7];

assign r_3 = r_2[9:7] + q_2[13] + q_3[18:13] + q_4[18:13] + q_5[18:13] + q_6[18:13] + q_7[18:13] + q_8[18:13] + q_9[18:13] + q_10[18:13] + q_11[18:13];

assign r_4 = r_3[9:7] + q_3[19] + q_4[24:19] + q_5[24:19] + q_6[24:19] + q_7[24:19] + q_8[24:19] + q_9[24:19] + q_10[24:19] + q_11[24:19];

assign r_5 = r_4[9:7] + q_4[25] + q_5[30:25] + q_6[30:25] + q_7[30:25] + q_8[30:25] + q_9[30:25] + q_10[30:25] + q_11[30:25];

assign r_6 = r_5[9:7] + q_5[31] + q_6[36:31] + q_7[36:31] + q_8[36:31] + q_9[36:31] + q_10[36:31] + q_11[36:31];

assign r_7 = r_6[8:7] + q_6[37] + q_7[42:37] + q_8[42:37] + q_9[42:37] + q_10[42:37] + q_11[42:37];

assign r_8 = r_7[8:7] + q_7[43] + q_8[48:43] + q_9[48:43] + q_10[48:43] + q_11[48:43];

assign r_9 = r_8[8:7] + q_8[49] + q_9[54:49] + q_10[54:49] + q_11[54:49];

assign r_10 = r_9[7] + q_9[55] + q_10[60:55] + q_11[60:55];

assign r_11 = r_10[7] + q_10[61] + q_11[63:61];


assign Q = {r_11, r_10[6:1], r_9[6:1], r_8[6:1], r_7[6:1], r_6[6:1], r_5[6:1], r_4[6:1], r_3[6:1], r_2[6:1], r_1[6:1]} + sum[6:3];


assign R = sum[2:1]; 

endmodule