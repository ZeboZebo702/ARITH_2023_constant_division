// Benchmark "q_10" written by ABC on Fri Jul 07 00:12:27 2023

module q_10 ( 
    x0, x1, x2, x3, x4,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64  );
  input  x0, x1, x2, x3, x4;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64;
  assign z00 = x0 & (x1 | (x2 & x3 & x4));
  assign z01 = x0 ? (~x1 & (~x2 | ~x3 | ~x4)) : (x1 & x2);
  assign z02 = x0 ? ((~x1 & (x2 ? ~x4 : x3)) | (x2 & (x4 ? (x1 | ~x3) : x3))) : (x1 ? ~x2 : (x2 & x3));
  assign z03 = (x2 & ((x0 & ~x4 & (x1 ^ x3)) | (~x1 & ~x3 & (~x0 | x4)))) | (~x0 & x4 & ((~x2 & x3) | (x1 & (~x2 | x3)))) | (~x2 & ((x1 & x3) | (x0 & ~x1 & ~x3)));
  assign z04 = (x2 & (x0 ? ((~x4 & (~x1 | ~x3)) | (x1 & x3 & x4)) : ((~x3 & x4) | (x1 & x3 & ~x4)))) | (~x2 & ((x4 & (~x0 ^ (~x1 | ~x3))) | (~x0 & ~x4 & (x1 ^ x3)))) | (x0 & ~x1 & ~x3 & ~x4);
  assign z05 = x3 ? ((x0 & (x1 ? x4 : (~x2 & ~x4))) | (~x0 & (x1 ? ~x4 : (x2 & x4))) | (x1 & (~x2 ^ ~x4))) : ((~x2 & (~x1 ^ ~x4)) | (~x1 & (x4 ? x0 : x2)));
  assign z06 = ((x0 | ~x3) & ((x2 & ~x4) | (x1 & ~x2 & x4))) | (~x0 & (x2 ? (x4 & (~x1 | x3)) : (x3 & ~x4))) | (~x3 & x4 & x0 & ~x2);
  assign z07 = ((x1 | ~x4) & (x0 ^ x3)) | (~x1 & x4 & (x0 ? (~x2 & x3) : ~x3));
  assign z08 = ~x1 ^ (~x4 | (x0 & x2 & x3));
  assign z09 = (x2 & (~x0 | ~x3 | ~x4)) | (x0 & x1 & ~x2 & x3 & x4);
  assign z10 = (x3 & (~x0 | ~x4 | (~x1 & ~x2))) | (~x3 & x4 & x0 & x1);
  assign z11 = (x4 & (~x0 | (~x1 & (~x2 | ~x3)))) | (x0 & x1 & ~x4);
  assign z60 = x1 ? ((x0 & ~x2 & (~x3 ^ x4)) | (x3 & ~x4 & (~x0 | x2))) : (x2 ? ((~x3 & ~x4) | (~x0 & x3 & x4)) : (~x3 & x4));
  assign z61 = x1 ? ((x0 & ~x2) ? (~x3 & x4) : (~x3 ^ x4)) : (x2 ? (~x3 & x4) : (x3 & ~x4));
  assign z12 = x0 ? (~x1 & (~x2 | ~x3 | ~x4)) : (x1 & x2);
  assign z13 = x0 ? ((~x1 & (x2 ? ~x4 : x3)) | (x2 & (x4 ? (x1 | ~x3) : x3))) : (x1 ? ~x2 : (x2 & x3));
  assign z14 = (x2 & ((x0 & ~x4 & (x1 ^ x3)) | (~x1 & ~x3 & (~x0 | x4)))) | (~x0 & x4 & ((~x2 & x3) | (x1 & (~x2 | x3)))) | (~x2 & ((x1 & x3) | (x0 & ~x1 & ~x3)));
  assign z15 = (x2 & (x0 ? ((~x4 & (~x1 | ~x3)) | (x1 & x3 & x4)) : ((~x3 & x4) | (x1 & x3 & ~x4)))) | (~x2 & ((x4 & (~x0 ^ (~x1 | ~x3))) | (~x0 & ~x4 & (x1 ^ x3)))) | (x0 & ~x1 & ~x3 & ~x4);
  assign z16 = x3 ? ((x0 & (x1 ? x4 : (~x2 & ~x4))) | (~x0 & (x1 ? ~x4 : (x2 & x4))) | (x1 & (~x2 ^ ~x4))) : ((~x2 & (~x1 ^ ~x4)) | (~x1 & (x4 ? x0 : x2)));
  assign z17 = ((x0 | ~x3) & ((x2 & ~x4) | (x1 & ~x2 & x4))) | (~x0 & (x2 ? (x4 & (~x1 | x3)) : (x3 & ~x4))) | (~x3 & x4 & x0 & ~x2);
  assign z18 = ((x1 | ~x4) & (x0 ^ x3)) | (~x1 & x4 & (x0 ? (~x2 & x3) : ~x3));
  assign z19 = ~x1 ^ (~x4 | (x0 & x2 & x3));
  assign z20 = (x2 & (~x0 | ~x3 | ~x4)) | (x0 & x1 & ~x2 & x3 & x4);
  assign z21 = (x3 & (~x0 | ~x4 | (~x1 & ~x2))) | (~x3 & x4 & x0 & x1);
  assign z22 = (x4 & (~x0 | (~x1 & (~x2 | ~x3)))) | (x0 & x1 & ~x4);
  assign z23 = x0 ? (~x1 & (~x2 | ~x3 | ~x4)) : (x1 & x2);
  assign z24 = x0 ? ((~x1 & (x2 ? ~x4 : x3)) | (x2 & (x4 ? (x1 | ~x3) : x3))) : (x1 ? ~x2 : (x2 & x3));
  assign z25 = (x2 & ((x0 & ~x4 & (x1 ^ x3)) | (~x1 & ~x3 & (~x0 | x4)))) | (~x0 & x4 & ((~x2 & x3) | (x1 & (~x2 | x3)))) | (~x2 & ((x1 & x3) | (x0 & ~x1 & ~x3)));
  assign z26 = (x2 & (x0 ? ((~x4 & (~x1 | ~x3)) | (x1 & x3 & x4)) : ((~x3 & x4) | (x1 & x3 & ~x4)))) | (~x2 & ((x4 & (~x0 ^ (~x1 | ~x3))) | (~x0 & ~x4 & (x1 ^ x3)))) | (x0 & ~x1 & ~x3 & ~x4);
  assign z27 = x3 ? ((x0 & (x1 ? x4 : (~x2 & ~x4))) | (~x0 & (x1 ? ~x4 : (x2 & x4))) | (x1 & (~x2 ^ ~x4))) : ((~x2 & (~x1 ^ ~x4)) | (~x1 & (x4 ? x0 : x2)));
  assign z28 = ((x0 | ~x3) & ((x2 & ~x4) | (x1 & ~x2 & x4))) | (~x0 & (x2 ? (x4 & (~x1 | x3)) : (x3 & ~x4))) | (~x3 & x4 & x0 & ~x2);
  assign z29 = ((x1 | ~x4) & (x0 ^ x3)) | (~x1 & x4 & (x0 ? (~x2 & x3) : ~x3));
  assign z30 = ~x1 ^ (~x4 | (x0 & x2 & x3));
  assign z31 = (x2 & (~x0 | ~x3 | ~x4)) | (x0 & x1 & ~x2 & x3 & x4);
  assign z32 = (x3 & (~x0 | ~x4 | (~x1 & ~x2))) | (~x3 & x4 & x0 & x1);
  assign z33 = (x4 & (~x0 | (~x1 & (~x2 | ~x3)))) | (x0 & x1 & ~x4);
  assign z34 = x0 ? (~x1 & (~x2 | ~x3 | ~x4)) : (x1 & x2);
  assign z35 = x0 ? ((~x1 & (x2 ? ~x4 : x3)) | (x2 & (x4 ? (x1 | ~x3) : x3))) : (x1 ? ~x2 : (x2 & x3));
  assign z36 = (x2 & ((x0 & ~x4 & (x1 ^ x3)) | (~x1 & ~x3 & (~x0 | x4)))) | (~x0 & x4 & ((~x2 & x3) | (x1 & (~x2 | x3)))) | (~x2 & ((x1 & x3) | (x0 & ~x1 & ~x3)));
  assign z37 = (x2 & (x0 ? ((~x4 & (~x1 | ~x3)) | (x1 & x3 & x4)) : ((~x3 & x4) | (x1 & x3 & ~x4)))) | (~x2 & ((x4 & (~x0 ^ (~x1 | ~x3))) | (~x0 & ~x4 & (x1 ^ x3)))) | (x0 & ~x1 & ~x3 & ~x4);
  assign z38 = x3 ? ((x0 & (x1 ? x4 : (~x2 & ~x4))) | (~x0 & (x1 ? ~x4 : (x2 & x4))) | (x1 & (~x2 ^ ~x4))) : ((~x2 & (~x1 ^ ~x4)) | (~x1 & (x4 ? x0 : x2)));
  assign z39 = ((x0 | ~x3) & ((x2 & ~x4) | (x1 & ~x2 & x4))) | (~x0 & (x2 ? (x4 & (~x1 | x3)) : (x3 & ~x4))) | (~x3 & x4 & x0 & ~x2);
  assign z40 = ((x1 | ~x4) & (x0 ^ x3)) | (~x1 & x4 & (x0 ? (~x2 & x3) : ~x3));
  assign z41 = ~x1 ^ (~x4 | (x0 & x2 & x3));
  assign z42 = (x2 & (~x0 | ~x3 | ~x4)) | (x0 & x1 & ~x2 & x3 & x4);
  assign z43 = (x3 & (~x0 | ~x4 | (~x1 & ~x2))) | (~x3 & x4 & x0 & x1);
  assign z44 = (x4 & (~x0 | (~x1 & (~x2 | ~x3)))) | (x0 & x1 & ~x4);
  assign z45 = x0 ? (~x1 & (~x2 | ~x3 | ~x4)) : (x1 & x2);
  assign z46 = x0 ? ((~x1 & (x2 ? ~x4 : x3)) | (x2 & (x4 ? (x1 | ~x3) : x3))) : (x1 ? ~x2 : (x2 & x3));
  assign z47 = (x2 & ((x0 & ~x4 & (x1 ^ x3)) | (~x1 & ~x3 & (~x0 | x4)))) | (~x0 & x4 & ((~x2 & x3) | (x1 & (~x2 | x3)))) | (~x2 & ((x1 & x3) | (x0 & ~x1 & ~x3)));
  assign z48 = (x2 & (x0 ? ((~x4 & (~x1 | ~x3)) | (x1 & x3 & x4)) : ((~x3 & x4) | (x1 & x3 & ~x4)))) | (~x2 & ((x4 & (~x0 ^ (~x1 | ~x3))) | (~x0 & ~x4 & (x1 ^ x3)))) | (x0 & ~x1 & ~x3 & ~x4);
  assign z49 = x3 ? ((x0 & (x1 ? x4 : (~x2 & ~x4))) | (~x0 & (x1 ? ~x4 : (x2 & x4))) | (x1 & (~x2 ^ ~x4))) : ((~x2 & (~x1 ^ ~x4)) | (~x1 & (x4 ? x0 : x2)));
  assign z50 = ((x0 | ~x3) & ((x2 & ~x4) | (x1 & ~x2 & x4))) | (~x0 & (x2 ? (x4 & (~x1 | x3)) : (x3 & ~x4))) | (~x3 & x4 & x0 & ~x2);
  assign z51 = ((x1 | ~x4) & (x0 ^ x3)) | (~x1 & x4 & (x0 ? (~x2 & x3) : ~x3));
  assign z52 = ~x1 ^ (~x4 | (x0 & x2 & x3));
  assign z53 = (x2 & (~x0 | ~x3 | ~x4)) | (x0 & x1 & ~x2 & x3 & x4);
  assign z54 = (x3 & (~x0 | ~x4 | (~x1 & ~x2))) | (~x3 & x4 & x0 & x1);
  assign z55 = (x4 & (~x0 | (~x1 & (~x2 | ~x3)))) | (x0 & x1 & ~x4);
  assign z56 = x0 ? (~x1 & (~x2 | ~x3 | ~x4)) : (x1 & x2);
  assign z57 = x0 ? ((~x1 & (x2 ? ~x4 : x3)) | (x2 & (x4 ? (x1 | ~x3) : x3))) : (x1 ? ~x2 : (x2 & x3));
  assign z58 = (x2 & ((x0 & ~x4 & (x1 ^ x3)) | (~x1 & ~x3 & (~x0 | x4)))) | (~x0 & x4 & ((~x2 & x3) | (x1 & (~x2 | x3)))) | (~x2 & ((x1 & x3) | (x0 & ~x1 & ~x3)));
  assign z59 = (x2 & (x0 ? ((~x4 & (~x1 | ~x3)) | (x1 & x3 & x4)) : ((~x3 & x4) | (x1 & x3 & ~x4)))) | (~x2 & ((x4 & (~x0 ^ (~x1 | ~x3))) | (~x0 & ~x4 & (x1 ^ x3)))) | (x0 & ~x1 & ~x3 & ~x4);
  assign z62 = x0 ? ((~x1 & (x2 ? ~x4 : x3)) | (x2 & (x4 ? (x1 | ~x3) : x3))) : (x1 ? ~x2 : (x2 & x3));
  assign z63 = (x2 & ((x0 & ~x4 & (x1 ^ x3)) | (~x1 & ~x3 & (~x0 | x4)))) | (~x0 & x4 & ((~x2 & x3) | (x1 & (~x2 | x3)))) | (~x2 & ((x1 & x3) | (x0 & ~x1 & ~x3)));
  assign z64 = (x2 & (x0 ? ((~x4 & (~x1 | ~x3)) | (x1 & x3 & x4)) : ((~x3 & x4) | (x1 & x3 & ~x4)))) | (~x2 & ((x4 & (~x0 ^ (~x1 | ~x3))) | (~x0 & ~x4 & (x1 ^ x3)))) | (x0 & ~x1 & ~x3 & ~x4);
endmodule


