// Benchmark "quot_res" written by ABC on Mon Feb 27 16:36:08 2023

module quot_res ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10;
  wire n24, n25, n26, n27, n28, n29, n30, n32, n33, n34, n35, n36, n37, n38,
    n39, n40, n41, n42, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
    n54, n55, n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82, n83,
    n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
    n98, n99, n100, n101, n102, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215;
  assign z00 = ~n27 | (x02 & (x03 | n24) & (~x03 | ~n25 | ~n26));
  assign n24 = x00 & ~x01;
  assign n25 = (~x00 | x01 | x04 | x05) & (x00 | ~x01 | ~x04 | ~x05);
  assign n26 = (~x00 | x01 | x04 | ~x05 | x06) & (x00 | ~x01 | ~x04 | x05 | ~x06);
  assign n27 = ~n30 & (x06 | ~n28 | ~n29 | (~x07 & ~x08));
  assign n28 = x03 & x02 & ~x00 & x01;
  assign n29 = x04 & ~x05;
  assign n30 = ~x02 & x00 & ~x01;
  assign z01 = n35 | n38 | n41 | (~x00 & ~n32);
  assign n32 = (x02 & x03 & x04 & (x01 | (~n33 & ~n34))) | (~x01 & (~x02 | ~x03 | (~x04 & ~n34)));
  assign n33 = x05 & x06;
  assign n34 = x07 & ~x06 & x04 & x05;
  assign n35 = n37 & ~n36 & x09 & ~x06 & ~x07;
  assign n36 = x00 ? (x04 | ~x08) : (~x04 | x08);
  assign n37 = x05 & x03 & ~x01 & x02;
  assign n38 = n40 & n39 & n24 & x02 & x03;
  assign n39 = ~x06 & x07;
  assign n40 = ~x04 & x05;
  assign n41 = n42 & (x01 ? (~x05 & ~x08) : (x05 & x08));
  assign n42 = ~x07 & ~x06 & x04 & x03 & ~x00 & x02;
  assign z02 = ~n55 | n53 | n50 | n44 | ~n49;
  assign n44 = n48 & (n45 | (~x06 & ~x08 & n40 & n47));
  assign n45 = n46 & ((x01 & ~x05 & (x02 ? (~x06 & ~x08) : (x06 & x08))) | (~x01 & ~x02 & x05 & x06 & x08));
  assign n46 = ~x00 & x04;
  assign n47 = x02 & x00 & ~x01;
  assign n48 = x03 & ~x07;
  assign n49 = (~x02 | ((x00 | (x03 & x04)) & (x01 | x03))) & (~x00 | x01 | x02 | ~x03 | ~x04);
  assign n50 = n52 & ~n51 & x06 & x07;
  assign n51 = (x00 | ~x04 | (~x01 ^ x05)) & (~x00 | x01 | x04 | ~x05);
  assign n52 = ~x02 & x03;
  assign n53 = ~n36 & n48 & n54 & (x02 ? (~x06 & ~x09) : (x06 & x09));
  assign n54 = ~x01 & x05;
  assign n55 = ~n56 & (n57 | ~n58 | ~x10 | ~n52);
  assign n56 = x03 & ((~x00 & x04 & (x01 ? (~x02 & x05) : (x02 & ~x05))) | (x00 & ~x01 & x02 & ~x04 & ~x05));
  assign n57 = (x00 | ~x04 | x08 | (x01 ? (x05 | ~x09) : (~x05 | x09))) & (~x00 | x01 | x04 | ~x05 | ~x08 | x09);
  assign n58 = x06 & ~x07;
  assign z03 = ~n60 | n66 | (~x07 & (n76 | (x05 & ~n72)));
  assign n60 = n63 & (x02 | n62) & (x03 | ~x07 | n61);
  assign n61 = (x01 | ((~x00 | ((~x02 | x04 | ~x05 | ~x06) & (x05 | x06 | x02 | ~x04))) & (x00 | ~x02 | ~x04 | ~x05 | ~x06))) & (x00 | ~x01 | ~x04 | (x02 ? (x05 | ~x06) : (~x05 | x06)));
  assign n62 = (x01 | ((~x00 | ((x03 | ~x04 | x05 | ~x06) & (~x05 | x06 | ~x03 | x04))) & (~x04 | ~x05 | x06 | x00 | ~x03))) & (x00 | ~x01 | ~x04 | (x03 ? (x05 | x06) : (~x05 | ~x06)));
  assign n63 = n65 & (n57 | ~n58 | (x10 ? ~n64 : ~n52));
  assign n64 = x02 & ~x03;
  assign n65 = (x01 | ((~x00 | x03 | ~x04 | (~x02 & ~x05)) & (~x03 | x05 | (x00 & x04)))) & (x00 | ((~x03 | x04) & (~x01 | ~x02 | x03 | ~x04 | ~x05)));
  assign n66 = ~x07 & (n70 | (~x01 & (n68 | (x05 & ~n67))));
  assign n67 = (~x00 | ~x03 | x04 | x08 | (~x02 ^ x06)) & (x00 | ~x02 | x03 | ~x04 | ~x06 | ~x08);
  assign n68 = n69 & n29 & x08 & x00 & ~x06;
  assign n69 = ~x02 & ~x03;
  assign n70 = n71 & ((x02 & ~x05 & (x03 ? (~x06 & ~x08) : (x06 & x08))) | (x05 & ~x06 & x08 & ~x02 & ~x03));
  assign n71 = x04 & ~x00 & x01;
  assign n72 = ~n74 & (~x04 | x06 | ~n73 | ~n69 | ~n75);
  assign n73 = ~x00 & x01;
  assign n74 = ~x01 & x02 & ~n36 & (x03 ? (~x06 & ~x09) : (x06 & x09));
  assign n75 = ~x08 & x09;
  assign n76 = n52 & n29 & n73 & ~x09 & x06 & ~x08;
  assign z04 = n82 | ~n85 | n98 | (~x07 & (~n78 | ~n90));
  assign n78 = (x04 | ~x06 | n81) & (x06 | (~n80 & (~x03 | n79)));
  assign n79 = (x04 | ((~x00 | x01 | (x02 ? (~x05 | x08) : (x05 | ~x08))) & (x00 | ~x01 | x02 | ~x05 | ~x08))) & (x00 | ~x01 | ~x02 | ~x04 | x05 | x08);
  assign n80 = n69 & ((~x04 & x08 & (x05 ? n73 : n24)) | (x04 & ~x05 & ~x08 & n24));
  assign n81 = (x01 | ~x05 | (x00 ? (x08 | (~x02 ^ x03)) : (~x02 | ~x08))) & (x00 | ~x01 | ~x02 | x05 | ~x08);
  assign n82 = ~x04 & ((~x03 & ~n84) | (~x00 & x02 & x03 & n83));
  assign n83 = x06 & x07 & (~x01 ^ ~x05);
  assign n84 = (x06 | (~x02 ^ x07) | (x00 ? (x01 | x05) : (~x01 | ~x05))) & (x00 | ~x02 | ~x06 | ~x07 | (~x01 ^ x05));
  assign n85 = ~n87 & ~n88 & ~n89 & ((x02 & x03) | n86 | (~x02 & ~x03));
  assign n86 = x00 ? (x01 | ((~x05 | (x04 ? (~x06 | ~x07) : x06)) & (x04 | (x06 ? x05 : ~x07)))) : ((~x01 | x04 | ~x05 | (~x06 & ~x07)) & (~x04 | ((x05 | x06) & (x01 | (x05 & x06)))));
  assign n87 = ~x01 & (x00 ? (~x04 & (x02 ? (x03 & ~x05) : (~x03 & x05))) : (x04 & (x02 ? (x03 & ~x05) : ~x03)));
  assign n88 = ~x00 & x01 & ((x02 & x03 & ~x04 & x05) | (~x02 & ~x03 & x04 & ~x05));
  assign n89 = ~x04 & x06 & n69 & (x00 ? (~x01 & ~x05) : (x01 & x05));
  assign n90 = x04 ? n91 : (~x05 | n94);
  assign n91 = x02 ? ((x03 | ~x06 | n92) & (x01 | ~x03 | ~n93)) : ((~x03 | ~x06 | n92) & (~x01 | x03 | ~n93));
  assign n92 = (x00 | ~x01 | x05 | x08 | x09) & (~x00 | x01 | ~x05 | ~x08 | ~x09);
  assign n93 = ~x09 & ~x08 & ~x06 & ~x00 & x05;
  assign n94 = (~n96 | ~n97) & (~x03 | x06 | ~n47 | ~n95);
  assign n95 = x08 & ~x09;
  assign n96 = x09 & (x01 ? (~x02 & ~x06) : (x02 & x06));
  assign n97 = ~x00 & ~x08;
  assign n98 = n58 & (n101 | ((~x02 | ~x03) & (x02 | x03) & (n99 | n100)));
  assign n99 = ~x09 & n54 & ((x00 & x08 & (~x04 ^ x10)) | (~x00 & x04 & ~x08 & ~x10));
  assign n100 = n71 & ~x10 & x09 & ~x05 & ~x08;
  assign n101 = ~n102 & x10 & ~x08 & ~x04 & ~x00 & x02;
  assign n102 = x01 ? (x05 | ~x09) : (~x05 | x09);
  assign z05 = (x03 & (~n114 | (~x07 & ~n104))) | ~n119 | (~x07 & ~n111);
  assign n104 = (n109 | ~n110) & (~n105 | n108 | (~n106 & ~n107));
  assign n105 = ~x05 & x06;
  assign n106 = x02 & ~x04;
  assign n107 = ~x02 & x04;
  assign n108 = (~x00 | x01 | ~x08 | ~x09) & (x08 | x09 | x00 | ~x01);
  assign n109 = (x00 | x08 | (x01 ? (x02 | x04) : (~x02 | ~x04))) & (~x00 | x01 | ~x02 | x04 | ~x08);
  assign n110 = ~x09 & x05 & ~x06;
  assign n111 = (~n97 | n112) & (~n24 | ~n105 | ~n113);
  assign n112 = (x05 | ((~x01 | ((x02 | x06 | ~x09) & (~x02 | x03 | ~x06 | x09))) & (x01 | ~x02 | ~x06 | ~x09))) & (~x01 | x02 | x03 | ~x05 | x06 | x09);
  assign n113 = x09 & x08 & x02 & ~x03;
  assign n114 = x01 ? (x00 | n118) : (~n115 & n116);
  assign n115 = x06 & ((x00 & ~x05 & x07 & (~x02 ^ ~x04)) | (~x00 & ~x02 & ~x04 & x05));
  assign n116 = (x04 | (x02 ? (~x05 | (~n117 & (x00 | x06))) : (x05 | ~n117))) & (x02 | ~x04 | ~x05 | ~n117);
  assign n117 = ~x08 & ~x07 & x00 & ~x06;
  assign n118 = (~x02 & (~x06 | (x05 & ~x07 & ~x08))) | (~x05 & (x04 | (x02 & ~x07 & ~x08))) | (x02 & x06 & (x07 | x08)) | (~x04 & x05) | (~x06 & ~x07 & ~x08);
  assign n119 = ~n122 & n126 & (x07 | (x02 & n120) | (~x02 & n121));
  assign n120 = (~x00 | x01 | x03 | ~x05 | ~x06 | x08) & (x00 | ((~x01 | ((~x05 | ~x06 | ~x08) & (x06 | x08 | ~x03 | x05))) & (x01 | x05 | ~x06 | ~x08)));
  assign n121 = (~x00 | x01 | ((~x05 | ((x06 | ~x08) & (~x03 | ~x06 | x08))) & (x03 | x05 | x06 | x08))) & (x00 | ~x01 | x05 | x06 | ~x08);
  assign n122 = n58 & ((~n123 & ~n124) | (~x01 & ~x09 & ~n125));
  assign n123 = (x00 | x08 | ((~x01 | ~x09 | (~x05 ^ ~x10)) & (x09 | x10 | x01 | ~x05))) & (~x00 | x01 | x05 | ~x08 | x09 | ~x10);
  assign n124 = x02 ^ (~x03 | ~x04);
  assign n125 = (x00 | ~x02 | x05 | x08 | ~x10) & (~x00 | ~x05 | ~x08 | x10 | (x02 ^ ~x03));
  assign n126 = ~n127 & (x03 | n128) & (~x05 | ~n30 | ~n39);
  assign n127 = ~x00 & ((x07 & ((x01 & (x02 ? (x05 & x06) : (~x05 & ~x06))) | (~x05 & x06 & ~x01 & x02))) | (~x01 & ~x02 & x05 & ~x06));
  assign n128 = ((~x02 ^ x06) | ((x01 | ~x05) & (x00 | ~x01 | x05))) & (~x00 | x01 | ~x02 | x05 | ~x06 | ~x07);
  assign z06 = ~n147 | (~x07 & (n138 | ~n140 | (~n130 & ~n131)));
  assign n130 = x06 ^ ~x10;
  assign n131 = ~n133 & (~x02 | n132) & (~x03 | (~n134 & ~n136));
  assign n132 = (x00 | x08 | (x03 & x04) | (~x01 ^ ~x09)) & (~x00 | x01 | x03 | ~x08 | x09);
  assign n133 = n95 & n30 & x03 & x04;
  assign n134 = n135 & ((x01 & ~x02 & x05 & x09) | (~x05 & ~x09 & ~x01 & x02));
  assign n135 = ~x08 & ~x00 & x04;
  assign n136 = n95 & n137 & n47;
  assign n137 = ~x04 & ~x05;
  assign n138 = ~n57 & n139;
  assign n139 = x03 & (x02 ? (~x06 & x10) : (x06 & ~x10));
  assign n140 = x03 ? (~n142 & n144 & (x06 | n141)) : n143;
  assign n141 = (x00 | x04 | x08 | (x01 ? (x02 | x09) : (~x02 | ~x09))) & (~x00 | x01 | x02 | ~x04 | ~x08 | ~x09);
  assign n142 = ~x04 & x06 & ~x08 & n73 & (~x02 ^ ~x09);
  assign n143 = (~x02 | ((x00 | x08 | (x01 ? (~x06 | x09) : (x06 | ~x09))) & (~x00 | x01 | x06 | ~x08 | ~x09))) & (x00 | ~x01 | x02 | x08 | (~x06 ^ ~x09));
  assign n144 = (x05 | x06 | ((~n106 | ~n145) & (~n135 | n146))) & (~x05 | ~x06 | ~n135 | n146);
  assign n145 = x09 & x08 & x00 & ~x01;
  assign n146 = x01 ? (x02 | x09) : (~x02 | ~x09);
  assign n147 = ~n148 & n157 & (x07 | (~n150 & ~n152 & n154));
  assign n148 = x03 & ((~x01 & ~n149) | (~x00 & x01 & ~x02 & n34));
  assign n149 = (x05 | ((x00 | x02 | ~x04 | ~x06) & (~x07 | ((~x00 | x04 | (~x02 ^ x06)) & (x00 | ~x02 | ~x04 | x06))))) & (x00 | ~x02 | ~x04 | ~x05 | ~x06 | ~x07);
  assign n150 = ~n151 & (~x02 ^ ~x08);
  assign n151 = (~x00 | x01 | ~x06 | (x03 & (x04 | x05))) & (x00 | ~x01 | ~x03 | ~x04 | ~x05 | x06);
  assign n152 = ~n153 & ((x03 & x04 & x06) | (~x06 & (~x03 | ~x04)));
  assign n153 = (~x00 | x01 | x02 | x08) & (x00 | ~x01 | ~x02 | ~x08);
  assign n154 = x06 ? ((~x05 | ~n156) & (~x01 | x02 | ~n155)) : ((x05 | ~n156) & (x01 | ~x02 | ~n155));
  assign n155 = ~x00 & x08 & (~x03 | ~x04);
  assign n156 = x08 & x04 & x03 & x02 & ~x00 & ~x01;
  assign n157 = x03 ? n159 : n158;
  assign n158 = (x00 | x01 | x02 | ~x06) & (~x07 | (x00 & x01) | (~x02 ^ x06));
  assign n159 = (x02 | ((x00 | x04 | ~x06 | (x01 & ~x07)) & (~x00 | x01 | ~x04 | x06 | ~x07))) & (x00 | ~x02 | ~x07 | ((~x01 | ~x04 | ~x06) & (x04 | x06)));
  assign z07 = n161 | n163 | ~n167 | ((x07 | ~x10) & ~n131 & (~x07 | x10));
  assign n161 = ~x03 & ((x04 & ~n162) | (~x04 & ~x07 & n47 & n75));
  assign n162 = (~x07 | ((x01 | ((~x00 | ~x08 | (~x02 ^ ~x09)) & (x08 | x09 | x00 | x02))) & (x00 | ~x01 | x02 | x08 | ~x09))) & (~x00 | x01 | ~x02 | x07 | x08);
  assign n163 = x03 & (n166 | (~x08 & (n165 | (n54 & ~n164))));
  assign n164 = (x00 | ~x04 | x09 | (x02 ? (~x06 | x07) : (x06 | ~x07))) & (~x00 | ~x02 | x04 | x06 | x07);
  assign n165 = x09 & n73 & n29 & (x02 ? n58 : n39);
  assign n166 = x08 & n24 & n39 & n40 & (~x02 ^ x09);
  assign n167 = n174 & ~n173 & ~n172 & ~n168 & n169;
  assign n168 = x03 & ~n57 & ((x07 & x10 & ~x02 & x06) | (~x07 & ~x10 & x02 & ~x06));
  assign n169 = (~x07 | ((~x08 | ~x09 | n170) & (x02 | x09 | n171))) & (x07 | x08 | x09 | n170);
  assign n170 = (~x00 | x01 | x04 | ~x05 | (x02 & x03)) & (x00 | ~x01 | ~x04 | x05);
  assign n171 = (x00 | ~x04 | x05 | (x01 ? ~x08 : (~x03 | x08))) & (~x00 | x01 | x03 | x04 | ~x05 | ~x08);
  assign n172 = n97 & (x01 ? (~x02 & ~x04 & (~x07 ^ x09)) : (x07 & x09 & (x02 | x04)));
  assign n173 = ~n25 & (x07 ? (x08 & (~x02 | x09)) : (~x08 & (~x09 | (x02 & x03))));
  assign n174 = (~x04 | (x07 ? (~x08 | n176) : (x08 | ~n30))) & ~n175 & (x04 | x07 | x08 | n176);
  assign n175 = ~x00 & x07 & ((~x04 & x08) | (~x01 & (x08 | (~x02 & ~x04))));
  assign n176 = (~x00 | x01 | x02 | ~x09) & (x00 | ~x01 | ~x02 | x09);
  assign z08 = n179 | ~n181 | n186 | n189 | (x02 & ~n178);
  assign n178 = (x01 | x09 | ((x00 | x08 | x10) & (x03 | (x00 ? (~x08 ^ x10) : (~x08 | ~x10))))) & (x00 | ~x01 | ~x09 | ((x08 | x10) & (x03 | ~x08 | ~x10)));
  assign n179 = n139 & (n180 | (~x05 & x07 & n71 & n75));
  assign n180 = ~x09 & n54 & ((~x00 & x04 & x07 & ~x08) | (x00 & ~x04 & (x07 ^ ~x08)));
  assign n181 = ~n182 & n184 & (~x03 | ~x08 | n183);
  assign n182 = ~x01 & (x00 ? (~x08 & ((~x03 & x09) | (~x02 & (~x03 | x09)))) : (x08 & (x09 | (~x02 & ~x03))));
  assign n183 = (~x00 | x01 | x02 | ~x04 | x09 | x10) & (x00 | x04 | (x01 ^ x09) | (~x02 ^ ~x10));
  assign n184 = (x09 | ((x00 | (x01 ? x08 : (~x08 | ~n185))) & (~x00 | x01 | x08 | ~n185))) & (x00 | ~x01 | ~x08 | ~x09 | (~n69 & ~n185));
  assign n185 = x10 & ~x02 & x03;
  assign n186 = x03 & (n188 | (~n187 & (~x02 ^ x10)));
  assign n187 = (x00 | ~x04 | ((x08 | ~x09 | ~x01 | ~x05) & (x01 | x05 | ~x08 | x09))) & (~x00 | x01 | x04 | x05 | x08 | x09);
  assign n188 = ~x05 & n24 & n106 & (x08 ? (~x09 & ~x10) : x09);
  assign n189 = x03 & (n190 | (~x06 & n24 & n40 & ~n191));
  assign n190 = n46 & ~n102 & ((x02 & x06 & ~x08 & x10) | (~x02 & ~x06 & x08 & ~x10));
  assign n191 = (~x02 | (x08 ? (x09 | x10) : ~x09)) & (x09 | x10 | x02 | x08);
  assign z09 = n193 | ~n197 | (~x01 & ~n196);
  assign n193 = x03 & ((n54 & ~n194) | (n73 & n29 & ~n195));
  assign n194 = (x06 | x10 | ((x00 | x02 | ~x04 | ~x09) & (~x00 | x04 | (~x02 ^ x09)))) & (x00 | ~x02 | ~x04 | ~x06 | x09 | ~x10);
  assign n195 = (x09 | x10 | x02 | x06) & (~x09 | ~x10 | ~x02 | ~x06);
  assign n196 = x09 ? (((x02 & ~x10) | (x03 & (x00 | x04))) & (x02 | ~x10)) : (x10 | ((~x00 | x02 | ~x03 | ~x04) & (~x02 | (x00 & x03))));
  assign n197 = ~n198 & ~n199 & (n203 | ~n204) & (~x03 | n201);
  assign n198 = n73 & ((~x09 & ((~x02 & x10) | ((~x03 | ~x04) & (~x02 | x10)))) | (x02 & x09 & ~x10));
  assign n199 = n200 & ((x00 & ~x01 & ~x04 & x05 & ~x09) | (~x00 & x04 & (x01 ? (~x05 & x09) : (x05 & ~x09))));
  assign n200 = x03 & x07 & (x02 ? (~x06 & x10) : (x06 & ~x10));
  assign n201 = (x09 | x10 | ~n137 | ~n47) & (~x09 | n202 | (x02 ^ x10));
  assign n202 = (~x00 | x01 | x04 | x05) & (x00 | ~x04 | (~x01 ^ ~x05));
  assign n203 = (~x00 | x01 | x04 | ~x05 | x08 | ~x09) & (x00 | ~x04 | ((~x01 | x05 | (~x08 ^ ~x09)) & (x01 | ~x05 | ~x08 | x09)));
  assign n204 = x03 & ~x07 & (x02 ? (~x06 & x10) : (x06 & ~x10));
  assign z10 = ~n211 | ~n213 | (n48 & (~n206 | n209 | n210));
  assign n206 = (~n54 | n207) & (~n73 | ~n29 | n208);
  assign n207 = x00 ? (x04 | x08 | (x02 ? (x06 | x10) : (~x06 | ~x10))) : (~x04 | ~x08 | (x02 ? (x06 | ~x10) : (~x06 | x10)));
  assign n208 = (x02 | ~x06 | ~x08 | x10) & (~x02 | x06 | (~x08 ^ ~x10));
  assign n209 = ~n36 & n54 & ((~x02 & x06 & x09 & ~x10) | (x02 & ~x06 & (x09 ^ ~x10)));
  assign n210 = n107 & n105 & n73 & x10 & ~x08 & ~x09;
  assign n211 = n212 & (n51 | ~n200);
  assign n212 = (~x00 | x01 | x02 | ~x03 | ~x04 | x10) & (((x00 | (x03 & x04)) & (x01 | x03)) | (~x02 ^ x10));
  assign n213 = ~x03 | (n214 & (~x10 | n215));
  assign n214 = (x01 | x05 | (~x02 ^ x10) | (x00 ^ ~x04)) & (x00 | ~x01 | ~x04 | ~x05 | (~x02 ^ ~x10));
  assign n215 = (x00 | ~x04 | (~x01 ^ x05) | (~x02 ^ ~x06)) & (~x00 | x01 | x02 | x04 | ~x05 | x06);
endmodule


