// Benchmark "q_3" written by ABC on Mon Feb 27 04:15:20 2023

module q_3 ( 
    x0, x1, x2, x3, x4, x5, x6,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28  );
  input  x0, x1, x2, x3, x4, x5, x6;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28;
  wire n38, n40, n41, n42, n44, n45, n47, n48, n50, n51, n52, n53, n54, n55,
    n56, n58, n59, n60, n61, n63, n64, n65, n67, n68, n70, n71, n72, n73,
    n74, n76, n78, n79, n80, n82, n83, n85, n86, n87, n89, n91, n92, n94,
    n95, n96, n97, n99, n100, n102, n103, n104, n105, n106, n107, n109,
    n110, n111, n112, n114, n115, n116, n117, n119, n120, n121, n122, n124,
    n125, n126, n127, n128, n130, n131, n132, n133, n134, n136, n137, n138,
    n139, n140, n141, n143, n144, n145, n146, n148, n149, n150, n151, n153,
    n154, n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166;
  assign z00 = x0 & x1 & x2 & ~n38;
  assign n38 = ~x6 & ~x5 & ~x3 & ~x4;
  assign z01 = ~n42 | (~x4 & n40 & n41);
  assign n40 = ~x5 & (x0 ? (~x3 & ~x6) : (x3 & x6));
  assign n41 = x1 & x2;
  assign n42 = x0 ? (x1 & x2) : (~x1 | ~x2 | ~x3 | (~x4 & ~x5));
  assign z02 = ~n45 | (n44 & (x1 ? (~x4 & ~x6) : (x4 & x6)));
  assign n44 = x2 & ~x5 & (x0 ^ x3);
  assign n45 = x1 ? (x2 & (x0 | x3)) : (~x2 | ((~x0 | (~x3 & (~x4 | ~x5))) & (~x3 | ~x4 | ~x5)));
  assign z03 = ~n48 | (n47 & (x2 ? (~x5 & ~x6) : (x5 & x6)));
  assign n47 = (x0 ^ x3) & (x1 ^ x4);
  assign n48 = x2 ? ((x0 | (x3 & (x1 | x4))) & (x1 | x3 | x4)) : ((~x0 | (~x3 & (~x1 | ~x4))) & (~x1 | ~x3 | ~x4));
  assign z04 = n50 | ~n51 | n55 | (~x6 & n47 & ~n56);
  assign n50 = (x1 ^ x4) & (x0 ? ((x3 & x5) | (~x2 & ~x3 & ~x5)) : (x2 ? (~x3 & x5) : (x3 & ~x5)));
  assign n51 = ~n52 & ~n53 & (~x0 | ~n41 | ~n54);
  assign n52 = x0 & (x1 ? (x3 & x4) : (~x3 & ~x4));
  assign n53 = ~x5 & x4 & x3 & x2 & x0 & ~x1;
  assign n54 = x6 & ~x5 & x3 & ~x4;
  assign n55 = ~x0 & (x1 ? (~x3 & x4) : (x3 & ~x4));
  assign n56 = ~x2 ^ x5;
  assign z05 = n59 | ~n60 | (x1 & ~n58);
  assign n58 = (x0 | ((x2 | ~x5 | (x3 ? x6 : (x4 | ~x6))) & (~x2 | x3 | x4 | x5 | ~x6))) & (~x3 | x6 | (x2 ? (x5 | (~x0 & x4)) : (~x4 | ~x5)));
  assign n59 = (x2 ^ x5) & (x1 ? ((x4 & x6) | (~x3 & ~x4 & ~x6)) : (x3 ? (~x4 & x6) : (x4 & ~x6)));
  assign n60 = x1 ? (x2 ? (~x4 | ~x5) : (x4 | x5)) : ((~x4 | ((x0 | n61 | (x2 & x5)) & (x2 | x5))) & (~x2 | x4 | ~x5));
  assign n61 = ~x3 ^ x6;
  assign z06 = ~n64 | (~n61 & ~n63);
  assign n63 = x2 ? (x5 ? ((~x1 | ~x4) & (~x0 | (~x1 & ~x4))) : ((x1 | x4) & (x0 | (x1 & x4)))) : ((~x5 | ((x1 | x4) & (x0 | (x1 & x4)))) & (~x0 | ~x4 | x5));
  assign n64 = x2 ? (x5 ? (~x6 | (~x3 & (x1 | n65))) : (x6 | (x3 & (~x1 | n65)))) : (x3 ? (x5 | ~x6) : (~x5 | x6));
  assign n65 = ~x0 ^ x4;
  assign z07 = (x3 & (x0 ? (x4 & x6) : (~x4 & ~x6))) | (~x3 & (x0 ? (x4 & ~x6) : (~x4 & x6))) | ((x0 ^ x4) & (~n67 | (x6 & n68)));
  assign n67 = (~x1 | ~x5 | (x3 ^ x6)) & (x1 | (x3 ? x6 : (x5 | ~x6))) & (~x3 | x5 | x6);
  assign n68 = (~x2 ^ x3) & (x1 ^ x5);
  assign z08 = (x0 & (x1 ? ((x4 & x5) | (~x2 & ~x4 & ~x5)) : (~x4 & (x2 ^ x5)))) | ~n70 | (~x0 & ((x4 & ((~x2 & ~x5) | (~x1 & (~x2 | ~x5)))) | (x1 & ~x4 & x5)));
  assign n70 = ~n71 & (~x0 | ~n72 | (~n73 & ~n74));
  assign n71 = (~x0 | (~x4 ^ x6)) & (x0 | (x4 ^ x6)) & x2 & (~x1 | ~x5) & (x1 | x5);
  assign n72 = ~x1 & ~x2;
  assign n73 = x6 & ~x4 & ~x5;
  assign n74 = ~x6 & ~x5 & x3 & ~x4;
  assign z09 = (~x1 & ((x2 & ~x5 & x6) | (x5 & (~x2 | ~x6)))) | (x1 & ((x2 & (~x5 ^ x6)) | (~x5 & (x6 ? ~x2 : x3)))) | (~x2 & ~x3 & ~x5 & ~x6 & ~n76);
  assign n76 = (~x1 | ~x4) & (~x0 | x1 | x4);
  assign z10 = ~n80 | ~n78 | (~x2 & n79 & ~x0 & x1);
  assign n78 = x6 ? x2 : (~x2 | (~x3 & ~x4));
  assign n79 = ~x6 & ~x5 & ~x3 & ~x4;
  assign n80 = x3 | x4 | x6 | ((~x2 | ~x5) & (~x0 | x2 | x5));
  assign z11 = n83 | ((x3 | (~x4 & (~x5 | n40))) & (x4 | x5 | n40 | ~n82));
  assign n82 = (x0 | x1 | ~x2 | x3 | x6) & (~x0 | ~x1 | x2 | ~x3 | ~x6);
  assign n83 = ~x4 & ~x5 & ((x0 & ~x1 & x3 & x6) | (~x0 & x1 & ~x3 & ~x6));
  assign z12 = n86 | ~n85 | (x3 & ~x4 & n87);
  assign n85 = (~x4 & (x5 | x6)) | (~x5 & ((x0 & x1 & x6) | (~x6 & (x4 | (~x0 & ~x1)))));
  assign n86 = ~x5 & ((x0 & x1 & ~x2 & x4 & x6) | (~x0 & ~x1 & x2 & ~x4 & ~x6));
  assign n87 = ~x5 & ((x0 & x1 & x2 & x6) | (~x0 & ~x1 & ~x2 & ~x6));
  assign z13 = ~n89 | (~x3 & x4 & n87);
  assign n89 = (~x0 & ((~x5 & x6) | (~x1 & ~x2 & ~x3 & ~x6))) | (x5 & (~x6 | (x0 & x1 & x2))) | (~x5 & x6 & (~x1 | ~x2 | ~x3));
  assign z14 = ~n92 | (~x3 & ~x4 & ~n91);
  assign n91 = (~x0 | ~x1 | ~x2 | (x5 ^ x6)) & (x0 | x1 | x2 | ~x5 | x6);
  assign n92 = (~x0 & (x6 | (~x1 & ~x2 & ~x3 & ~x4))) | (x6 & (~x1 | ~x2 | (~x3 & ~x4))) | (x0 & x1 & x2 & ~x6);
  assign z15 = ~n94 | ((x1 | (~x0 & (x2 | x3 | x4))) & (~x0 | (x2 & (x3 | x4))) & (~x2 | ~x3 | x0 | ~x1));
  assign n94 = ~n96 & (x5 | ~n95 | n97);
  assign n95 = ~x0 & ~x4;
  assign n96 = ~x3 & ~x4 & x5 & (x0 ? (x1 & x2) : (~x1 & ~x2));
  assign n97 = (~x1 | ~x2 | ~x3 | x6) & (x1 | x2 | x3 | ~x6);
  assign z16 = ~n100 | (~x5 & ~n99);
  assign n99 = (x0 | ((x1 | ((x2 | x3 | x4 | ~x6) & (~x2 | ~x3 | ~x4 | x6))) & (~x1 | ~x2 | ~x3 | x4 | ~x6))) & (~x0 | x1 | ~x2 | x3 | ~x4 | x6);
  assign n100 = (~x1 & x2 & ((x3 & x4) | (x0 & (x3 | x4)))) | (~x2 & (x1 | (~x4 & ~x5 & ~x0 & ~x3))) | (x1 & ((~x3 & ~x4 & ~x5) | (~x0 & (~x3 | (~x4 & ~x5)))));
  assign z17 = ~n102 | ~n103 | ~n105;
  assign n102 = (x1 | x2 | (x0 ? (x3 | x4) : (~x3 ^ x4))) & (~x0 | ~x1 | ~x2 | (~x3 & ~x4));
  assign n103 = x2 ? (~x5 | ~n47) : ((x5 | ~n47) & (x3 | x4 | n104));
  assign n104 = (~x0 | ~x1 | ~x5 | x6) & (x0 | x1 | x5 | ~x6);
  assign n105 = n107 & (n106 | (x2 ? (x5 | ~x6) : (~x5 | x6)));
  assign n106 = (x0 | ~x3 | (~x1 ^ x4)) & (~x0 | x1 | x3 | ~x4);
  assign n107 = (x0 | ((x2 | x3 | x4 | ~x5) & (~x1 | (x2 ? (~x3 | ~x4) : x3)))) & (~x2 | ~x3 | ~x0 | x1);
  assign z18 = n110 | ~n111 | (~x4 & ~n109) | ~n112;
  assign n109 = (~x1 | (x0 ? ((~x5 | ~x6 | x2 | x3) & (x5 | x6 | ~x2 | ~x3)) : (~x3 | ~x6 | (~x2 ^ x5)))) & (x3 | x5 | ~x6 | x0 | x1 | x2);
  assign n110 = (x0 | ((~x2 | x3 | ~x5) & (~x3 | x5))) & (~x5 | ((x2 | ~x3) & (~x0 | (x2 & ~x3)))) & (~x1 | ~x4) & (x1 | x4) & (x5 | (x3 ? ~x2 : ~x0));
  assign n111 = x0 | (x1 ? (~x3 | ~x4) : (x3 | x4 | (~x2 & ~x5)));
  assign n112 = (x1 | ~x3 | ((~x0 | x4) & (x0 | ~x4 | ~x6 | n56))) & (~x0 | x3 | ~x4 | (~x1 & (~x6 | n56)));
  assign z19 = n115 | ~n116 | (~x5 & ~n114) | ~n117;
  assign n114 = (x1 | ((~x0 | ~x2 | ~x4 | (~x3 ^ x6)) & (x3 | x4 | ~x6 | x0 | x2))) & (x0 | ~x1 | ~x2 | ~x3 | ~x4 | x6);
  assign n115 = (x1 | ((~x3 | x4 | ~x6) & (~x4 | x6))) & (~x6 | ((x3 | ~x4) & (~x1 | (x3 & ~x4)))) & (~x2 | ~x5) & (x2 | x5) & (x6 | (x4 ? ~x3 : ~x1));
  assign n116 = x1 | (x2 ? (~x4 | ~x5) : (x4 | x5 | (~x0 & ~x3)));
  assign n117 = (~x5 | ((~x0 | n61 | (x1 ? x4 : (x2 | ~x4))) & (~x1 | ~x2 | x4))) & (~x1 | x2 | ~x4 | x5);
  assign z20 = (~x6 & (~n119 | (x3 & ~n120))) | ~n121 | (~x3 & x6 & ~n120);
  assign n119 = (~x0 | ((x2 | x3 | x5) & (~x3 | x4 | ~x5 | x1 | ~x2))) & (x2 | x3 | x5 | (~x1 & ~x4)) & (~x3 | ~x4 | ~x5 | x0 | x1 | ~x2);
  assign n120 = (x0 | (x2 ? (x4 | ~x5) : x5)) & (x2 | (x5 ? ((~x1 | ~x4) & (~x0 | (~x1 & ~x4))) : x4)) & (~x4 | x5 | ~x0 | ~x2);
  assign n121 = (~x2 | (x3 ? (x5 | ~x6) : (~x5 | x6))) & (~x6 | ((x2 | ~x3 | ~x5) & (x5 | ~n122 | x3 | ~x4)));
  assign n122 = x2 & ~x0 & x1;
  assign z21 = n125 | n126 | n127 | n128 | (x6 & ~n124);
  assign n124 = (~x3 & (~x2 | (~x4 & ~x5))) | (~x0 & ~x4) | (~x1 & ~x5) | (x2 & x3) | (x0 & x4) | (x1 & x5);
  assign n125 = (~x1 | ((x5 | ~x6) & (x3 | ~x5 | x6))) & (x1 | (x6 ? ~x5 : ~x3)) & (~x3 | (~x5 ^ ~x6)) & (x3 | x5 | ~x6) & (x0 | x4) & (~x0 | ~x4);
  assign n126 = ~x1 & ~x2 & ((x0 & x4 & (x3 ^ x6)) | (~x4 & x6 & ~x0 & x3));
  assign n127 = (~x3 | (~x4 ^ ~x6)) & (x3 | (~x4 ^ x6)) & (~x0 | x4) & (x1 | x2) & (x0 | ~x4);
  assign n128 = n72 & ~x6 & x5 & ~x4 & ~x0 & ~x3;
  assign z22 = n131 | n133 | (~x3 & ~n130) | ~n134;
  assign n130 = x1 ? (~x2 | x5 | (x0 ? (~x4 | x6) : (x4 ^ x6))) : ((~x5 | ((~x0 | ~x4 | (x2 ^ ~x6)) & (x0 | ~x2 | x4 | x6))) & (x4 | ~x6 | x0 | x2));
  assign n131 = ~n132 & (x1 ? (x3 & ~x5) : x5);
  assign n132 = x0 ? (x2 ? (x4 | ~x6) : (~x4 | x6)) : (x2 ? (~x4 | ~x6) : (x4 | x6));
  assign n133 = ~x2 & ~x5 & ((~x0 & ~x4 & (x1 ^ x3)) | (x0 & x1 & ~x3 & x4));
  assign n134 = x0 ? (x1 ? (x4 | ~x5) : (~x4 | x5)) : ((~x1 | ((~x4 | ~x5) & (~x2 | ~n74))) & (x4 | x5 | x1 | ~x2));
  assign z23 = n137 | ~n138 | ~n139 | ((~x4 | ~x6) & ~n136 & (x4 | x6));
  assign n136 = (x1 | x2 | x3 | x5) & (~x1 | ~x3 | (x0 ? (~x2 | x5) : (x2 | ~x5)));
  assign n137 = ~x5 & n72 & ((~x0 & x4 & (x3 ^ x6)) | (x0 & x3 & ~x4 & x6));
  assign n138 = x1 ? ((x0 | ~x2 | ~x4 | x5 | ~x6) & (~x0 | x2 | x4 | ~x5 | x6)) : (x0 ? (x4 | ((x5 | x6) & (~x2 | ~x5 | ~x6))) : (~x2 | ~x4 | (~x5 ^ ~x6)));
  assign n139 = (n140 | (~x0 ^ ~x4)) & (~x1 | ~x5 | n141);
  assign n140 = (x1 & ((x2 & (x6 ? x5 : x3)) | (~x5 & ~x6) | (x3 & x5 & x6))) | (~x1 & ((~x2 & (~x3 | (x5 & ~x6))) | (~x5 & x6) | (~x3 & x5 & ~x6))) | (~x5 & (x2 ? (x3 & ~x6) : ~x3));
  assign n141 = (x3 | ((~x0 | x4 | (~x2 ^ x6)) & (x0 | x2 | ~x4 | x6))) & (x0 | ~x2 | ~x3 | x4 | x6);
  assign z24 = n144 | n145 | (x2 ? ~n146 : ~n143);
  assign n143 = (((x0 | ~x3 | (~x1 ^ x4)) & (~x0 | x1 | x3 | ~x4)) | (~x5 ^ x6)) & (~x1 | (~x5 ^ ~x6) | (x0 ? (~x3 | x4) : ~x4)) & (x0 | x1 | x3 | x4 | ~x5 | x6);
  assign n144 = ~x4 & ((x1 & ((~x2 & ~x3 & ~x6) | (~x0 & x2 & x6))) | (~x0 & ((x2 & ~x3 & x6) | (~x1 & x3 & (~x2 ^ ~x6)))) | (x0 & ~x1 & ~x2 & ~x6));
  assign n145 = x4 & ((x0 & (x2 ? (x3 ^ x6) : ((x3 & x6) | (x1 & ~x3 & ~x6)))) | (~x0 & ~x1 & ~x2 & ~x3 & ~x6));
  assign n146 = (~x4 | ((x0 | (x1 ? (~x5 | x6) : (x5 | ~x6))) & (~x0 | ~x1 | ~x3 | ~x5 | ~x6))) & (~x0 | x4 | (x1 ? (~x5 | (x3 ^ ~x6)) : (x5 | ~x6)));
  assign z25 = n55 | n149 | ~n150 | ~n151 | (x6 & ~n148);
  assign n148 = x1 ? ((x3 | x4 | ~x5 | x0 | x2) & (~x2 | ((x0 | (x3 ? (~x4 | ~x5) : (x4 | x5))) & (~x0 | ~x3 | ~x4 | x5)))) : (x0 ? (~x3 | (x2 ? (x4 | ~x5) : (~x4 | x5))) : (x3 | ~x4 | (x2 ^ ~x5)));
  assign n149 = (~x0 | ((x3 | ~x5) & (x2 | ~x3 | x5))) & (x5 | ((~x2 | x3) & (x0 | (~x2 & x3)))) & (~x1 | ~x4) & (x1 | x4) & (~x5 | (x3 ? x0 : x2));
  assign n150 = ~x0 | ((x1 | x3 | x4) & (~x3 | ~x4 | ~x1 | x2));
  assign n151 = ~x0 | x6 | ~n41 | (x3 ? ~x4 : (x4 | x5));
  assign z26 = ~n155 | (x0 ? ~n153 : ~n154);
  assign n153 = (~x3 | ((~x4 | (x1 ? (x2 ? (~x5 | x6) : (x5 | ~x6)) : (x2 ? (~x5 | ~x6) : (x5 | x6)))) & (x1 | ~x2 | x4 | ~x5 | x6))) & (x1 | x3 | x4 | ~x6 | (~x2 ^ x5));
  assign n154 = (x3 | (x4 ? ((~x1 | ~x2 | x5 | ~x6) & (x1 | x2 | ~x5 | x6)) : ((~x2 ^ x5) | (x1 ^ ~x6)))) & (~x1 | ~x2 | ~x3 | ~x4 | ~x5 | x6);
  assign n155 = ~n156 & ~n158 & (n157 | (x0 ? (~x1 | x4) : (x1 | ~x4)));
  assign n156 = ~x0 & (x1 ? ((~x2 & (x4 ^ ~x5)) | (x4 & ((~x3 & x5) | (x2 & x3 & ~x5)))) : (~x4 & ((x3 & x5) | (x2 & (x3 | x5)))));
  assign n157 = (x5 | (x2 & (x3 | x6))) & (~x2 | ~x3 | ~x5 | ~x6);
  assign n158 = x0 & (((~x2 ^ ~x5) & (x1 ? x4 : (x3 & ~x4))) | (~x3 & (x1 ? (x4 & x5) : (x2 ? (~x4 & x5) : (x4 & ~x5)))));
  assign z27 = n161 | ~n163 | n165 | n166 | (x2 & ~n160);
  assign n160 = (~x0 | ((~x1 | ~x3 | x4 | x5 | ~x6) & (x1 | x3 | ~x4 | ~x5 | x6))) & (x3 | ~x4 | x6 | x0 | ~x1);
  assign n161 = ~n162 & (x3 ? (x4 & x6) : (~x4 & ~x6));
  assign n162 = (x5 & ((x0 & x1) | x2)) | (~x0 & ~x1) | (~x2 & ~x5);
  assign n163 = ((~x3 ^ x6) | (~x2 ^ ~x5)) & (~x2 | ((~x5 | ~x6 | ~n95) & (x3 | x6 | n164))) & (~x6 | n164 | x2 | ~x3);
  assign n164 = x0 ? (~x1 | ~x5) : (x1 | x5);
  assign n165 = ~x0 & ~x2 & ((x1 & x3 & ~x5 & x6) | (~x1 & ~x3 & x5 & ~x6));
  assign n166 = x0 & ~x2 & ~x5 & (x3 ? (~x4 & x6) : (x4 & ~x6));
  assign z28 = n125 | n126 | n127 | n128 | (x6 & ~n124);
endmodule


