module div_16_3(X, Q, R );

input  [16:1] X;
output [15:1] Q;  
output [2:1] R;  

//wire [28:1] Q_temp;

wire [8:1] r_1;
wire [7:1] r_2;
wire [3:1] r_3;

wire [4:1] sum_res;
wire [4:1] sum;

wire [9:1] q_1;
wire [15:1] q_2;
wire [17:1] q_3;


q_1 label1 ( .x0(X[8]),.x1(X[7]),.x2(X[6]),.x3(X[5]),.x4(X[4]),.x5(X[3]),
.z0(q_1[9]),.z1(q_1[8]),.z2(q_1[7]),.z3(q_1[6]),.z4(q_1[5]),.z5(q_1[4]),.z6(q_1[3]),.z7(q_1[2]),.z8(q_1[1]));

q_2 label2 ( .x0(X[14]),.x1(X[13]),.x2(X[12]),.x3(X[11]),.x4(X[10]),.x5(X[9]),
.z00(q_2[15]),.z01(q_2[14]),.z02(q_2[13]),.z03(q_2[12]),.z04(q_2[11]),.z05(q_2[10]),.z06(q_2[9]),.z07(q_2[8]),.z08(q_2[7]),.z09(q_2[6]),.z10(q_2[5]),.z11(q_2[4]),.z12(q_2[3]),.z13(q_2[2]),.z14(q_2[1]));

q_3 label3 ( .x0(X[16]),.x1(X[15]),
.z00(q_3[17]),.z01(q_3[16]),.z02(q_3[15]),.z03(q_3[14]),.z04(q_3[13]),.z05(q_3[12]),.z06(q_3[11]),.z07(q_3[10]),.z08(q_3[9]),.z09(q_3[8]),.z10(q_3[7]),.z11(q_3[6]),.z12(q_3[5]),.z13(q_3[4]),.z14(q_3[3]),.z15(q_3[2]),.z16(q_3[1]));


assign sum_res = X[2:1] + q_1[2:1] + q_2[2:1] + q_3[2:1];

quot_res  label10 (.x0(sum_res[4]),.x1(sum_res[3]),.x2(sum_res[2]),.x3(sum_res[1]),
                  .z0(sum[4]),.z1(sum[3]),.z2(sum[2]),.z3(sum[1]));


assign r_1 = q_1[8:3] + q_2[8:3] + q_3[8:3];

assign r_2 = r_1[8:7] + q_1[9] + q_2[14:9] + q_3[14:9];

assign r_3 = r_2[7] + q_2[15] + q_3[17:15];


assign Q = {r_3, r_2[6:1], r_1[6:1]} + sum[4:3];


//assign Q = Q_temp;

assign R = sum[2:1]; 

endmodule