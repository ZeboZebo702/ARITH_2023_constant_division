module div_64_5(X, Q, R );

input  [64:1] X;
output [62:1] Q;  
output [3:1] R;  


wire [10:1] r_1;
wire [9:1] r_2;
wire [9:1] r_3;
wire [9:1] r_4;
wire [9:1] r_5;
wire [9:1] r_6;
wire [8:1] r_7;
wire [8:1] r_8;
wire [8:1] r_9;
wire [7:1] r_10;
wire [2:1] r_11;


wire [6:1] sum_res;
wire [7:1] sum;

wire [10:1] q_1;
wire [16:1] q_2;
wire [22:1] q_3;
wire [28:1] q_4;
wire [34:1] q_5;
wire [40:1] q_6;
wire [46:1] q_7;
wire [52:1] q_8;
wire [58:1] q_9;
wire [64:1] q_10;
wire [64:1] q_11;


q_1 label1 ( .x0(X[9]),.x1(X[8]),.x2(X[7]),.x3(X[6]),.x4(X[5]),.x5(X[4]),
.z0(q_1[10]),.z1(q_1[9]),.z2(q_1[8]),.z3(q_1[7]),.z4(q_1[6]),.z5(q_1[5]),.z6(q_1[4]),.z7(q_1[3]),.z8(q_1[2]),.z9(q_1[1]));

q_2 label2 ( .x0(X[15]),.x1(X[14]),.x2(X[13]),.x3(X[12]),.x4(X[11]),.x5(X[10]),
.z00(q_2[16]),.z01(q_2[15]),.z02(q_2[14]),.z03(q_2[13]),.z04(q_2[12]),.z05(q_2[11]),.z06(q_2[10]),.z07(q_2[9]),.z08(q_2[8]),.z09(q_2[7]),.z10(q_2[6]),.z11(q_2[5]),.z12(q_2[4]),.z13(q_2[3]),.z14(q_2[2]),.z15(q_2[1]));

q_3 label3 ( .x0(X[21]),.x1(X[20]),.x2(X[19]),.x3(X[18]),.x4(X[17]),.x5(X[16]),
.z00(q_3[22]),.z01(q_3[21]),.z02(q_3[20]),.z03(q_3[19]),.z04(q_3[18]),.z05(q_3[17]),.z06(q_3[16]),.z07(q_3[15]),.z08(q_3[14]),.z09(q_3[13]),.z10(q_3[12]),.z11(q_3[11]),.z12(q_3[10]),.z13(q_3[9]),.z14(q_3[8]),.z15(q_3[7]),.z16(q_3[6]),.z17(q_3[5]),.z18(q_3[4]),.z19(q_3[3]),.z20(q_3[2]),.z21(q_3[1]));

q_4 label4 ( .x0(X[27]),.x1(X[26]),.x2(X[25]),.x3(X[24]),.x4(X[23]),.x5(X[22]),
.z00(q_4[28]),.z01(q_4[27]),.z02(q_4[26]),.z03(q_4[25]),.z04(q_4[24]),.z05(q_4[23]),.z06(q_4[22]),.z07(q_4[21]),.z08(q_4[20]),.z09(q_4[19]),.z10(q_4[18]),.z11(q_4[17]),.z12(q_4[16]),.z13(q_4[15]),.z14(q_4[14]),.z15(q_4[13]),.z16(q_4[12]),.z17(q_4[11]),.z18(q_4[10]),.z19(q_4[9]),.z20(q_4[8]),.z21(q_4[7]),.z22(q_4[6]),.z23(q_4[5]),.z24(q_4[4]),.z25(q_4[3]),.z26(q_4[2]),.z27(q_4[1]));

q_5 label5 ( .x0(X[33]),.x1(X[32]),.x2(X[31]),.x3(X[30]),.x4(X[29]),.x5(X[28]),
.z00(q_5[34]),.z01(q_5[33]),.z02(q_5[32]),.z03(q_5[31]),.z04(q_5[30]),.z05(q_5[29]),.z06(q_5[28]),.z07(q_5[27]),.z08(q_5[26]),.z09(q_5[25]),.z10(q_5[24]),.z11(q_5[23]),.z12(q_5[22]),.z13(q_5[21]),.z14(q_5[20]),.z15(q_5[19]),.z16(q_5[18]),.z17(q_5[17]),.z18(q_5[16]),.z19(q_5[15]),.z20(q_5[14]),.z21(q_5[13]),.z22(q_5[12]),.z23(q_5[11]),.z24(q_5[10]),.z25(q_5[9]),.z26(q_5[8]),.z27(q_5[7]),.z28(q_5[6]),.z29(q_5[5]),.z30(q_5[4]),.z31(q_5[3]),.z32(q_5[2]),.z33(q_5[1]));

q_6 label6 ( .x0(X[39]),.x1(X[38]),.x2(X[37]),.x3(X[36]),.x4(X[35]),.x5(X[34]),
.z00(q_6[40]),.z01(q_6[39]),.z02(q_6[38]),.z03(q_6[37]),.z04(q_6[36]),.z05(q_6[35]),.z06(q_6[34]),.z07(q_6[33]),.z08(q_6[32]),.z09(q_6[31]),.z10(q_6[30]),.z11(q_6[29]),.z12(q_6[28]),.z13(q_6[27]),.z14(q_6[26]),.z15(q_6[25]),.z16(q_6[24]),.z17(q_6[23]),.z18(q_6[22]),.z19(q_6[21]),.z20(q_6[20]),.z21(q_6[19]),.z22(q_6[18]),.z23(q_6[17]),.z24(q_6[16]),.z25(q_6[15]),.z26(q_6[14]),.z27(q_6[13]),.z28(q_6[12]),.z29(q_6[11]),.z30(q_6[10]),.z31(q_6[9]),.z32(q_6[8]),.z33(q_6[7]),.z34(q_6[6]),.z35(q_6[5]),.z36(q_6[4]),.z37(q_6[3]),.z38(q_6[2]),.z39(q_6[1]));

q_7 label7 ( .x0(X[45]),.x1(X[44]),.x2(X[43]),.x3(X[42]),.x4(X[41]),.x5(X[40]),
.z00(q_7[46]),.z01(q_7[45]),.z02(q_7[44]),.z03(q_7[43]),.z04(q_7[42]),.z05(q_7[41]),.z06(q_7[40]),.z07(q_7[39]),.z08(q_7[38]),.z09(q_7[37]),.z10(q_7[36]),.z11(q_7[35]),.z12(q_7[34]),.z13(q_7[33]),.z14(q_7[32]),.z15(q_7[31]),.z16(q_7[30]),.z17(q_7[29]),.z18(q_7[28]),.z19(q_7[27]),.z20(q_7[26]),.z21(q_7[25]),.z22(q_7[24]),.z23(q_7[23]),.z24(q_7[22]),.z25(q_7[21]),.z26(q_7[20]),.z27(q_7[19]),.z28(q_7[18]),.z29(q_7[17]),.z30(q_7[16]),.z31(q_7[15]),.z32(q_7[14]),.z33(q_7[13]),.z34(q_7[12]),.z35(q_7[11]),.z36(q_7[10]),.z37(q_7[9]),.z38(q_7[8]),.z39(q_7[7]),.z40(q_7[6]),.z41(q_7[5]),.z42(q_7[4]),.z43(q_7[3]),.z44(q_7[2]),.z45(q_7[1]));

q_8 label8 ( .x0(X[51]),.x1(X[50]),.x2(X[49]),.x3(X[48]),.x4(X[47]),.x5(X[46]),
.z00(q_8[52]),.z01(q_8[51]),.z02(q_8[50]),.z03(q_8[49]),.z04(q_8[48]),.z05(q_8[47]),.z06(q_8[46]),.z07(q_8[45]),.z08(q_8[44]),.z09(q_8[43]),.z10(q_8[42]),.z11(q_8[41]),.z12(q_8[40]),.z13(q_8[39]),.z14(q_8[38]),.z15(q_8[37]),.z16(q_8[36]),.z17(q_8[35]),.z18(q_8[34]),.z19(q_8[33]),.z20(q_8[32]),.z21(q_8[31]),.z22(q_8[30]),.z23(q_8[29]),.z24(q_8[28]),.z25(q_8[27]),.z26(q_8[26]),.z27(q_8[25]),.z28(q_8[24]),.z29(q_8[23]),.z30(q_8[22]),.z31(q_8[21]),.z32(q_8[20]),.z33(q_8[19]),.z34(q_8[18]),.z35(q_8[17]),.z36(q_8[16]),.z37(q_8[15]),.z38(q_8[14]),.z39(q_8[13]),.z40(q_8[12]),.z41(q_8[11]),.z42(q_8[10]),.z43(q_8[9]),.z44(q_8[8]),.z45(q_8[7]),.z46(q_8[6]),.z47(q_8[5]),.z48(q_8[4]),.z49(q_8[3]),.z50(q_8[2]),.z51(q_8[1]));

q_9 label9 ( .x0(X[57]),.x1(X[56]),.x2(X[55]),.x3(X[54]),.x4(X[53]),.x5(X[52]),
.z00(q_9[58]),.z01(q_9[57]),.z02(q_9[56]),.z03(q_9[55]),.z04(q_9[54]),.z05(q_9[53]),.z06(q_9[52]),.z07(q_9[51]),.z08(q_9[50]),.z09(q_9[49]),.z10(q_9[48]),.z11(q_9[47]),.z12(q_9[46]),.z13(q_9[45]),.z14(q_9[44]),.z15(q_9[43]),.z16(q_9[42]),.z17(q_9[41]),.z18(q_9[40]),.z19(q_9[39]),.z20(q_9[38]),.z21(q_9[37]),.z22(q_9[36]),.z23(q_9[35]),.z24(q_9[34]),.z25(q_9[33]),.z26(q_9[32]),.z27(q_9[31]),.z28(q_9[30]),.z29(q_9[29]),.z30(q_9[28]),.z31(q_9[27]),.z32(q_9[26]),.z33(q_9[25]),.z34(q_9[24]),.z35(q_9[23]),.z36(q_9[22]),.z37(q_9[21]),.z38(q_9[20]),.z39(q_9[19]),.z40(q_9[18]),.z41(q_9[17]),.z42(q_9[16]),.z43(q_9[15]),.z44(q_9[14]),.z45(q_9[13]),.z46(q_9[12]),.z47(q_9[11]),.z48(q_9[10]),.z49(q_9[9]),.z50(q_9[8]),.z51(q_9[7]),.z52(q_9[6]),.z53(q_9[5]),.z54(q_9[4]),.z55(q_9[3]),.z56(q_9[2]),.z57(q_9[1]));

q_10 label10 ( .x0(X[63]),.x1(X[62]),.x2(X[61]),.x3(X[60]),.x4(X[59]),.x5(X[58]),
.z00(q_10[64]),.z01(q_10[63]),.z02(q_10[62]),.z03(q_10[61]),.z04(q_10[60]),.z05(q_10[59]),.z06(q_10[58]),.z07(q_10[57]),.z08(q_10[56]),.z09(q_10[55]),.z10(q_10[54]),.z11(q_10[53]),.z12(q_10[52]),.z13(q_10[51]),.z14(q_10[50]),.z15(q_10[49]),.z16(q_10[48]),.z17(q_10[47]),.z18(q_10[46]),.z19(q_10[45]),.z20(q_10[44]),.z21(q_10[43]),.z22(q_10[42]),.z23(q_10[41]),.z24(q_10[40]),.z25(q_10[39]),.z26(q_10[38]),.z27(q_10[37]),.z28(q_10[36]),.z29(q_10[35]),.z30(q_10[34]),.z31(q_10[33]),.z32(q_10[32]),.z33(q_10[31]),.z34(q_10[30]),.z35(q_10[29]),.z36(q_10[28]),.z37(q_10[27]),.z38(q_10[26]),.z39(q_10[25]),.z40(q_10[24]),.z41(q_10[23]),.z42(q_10[22]),.z43(q_10[21]),.z44(q_10[20]),.z45(q_10[19]),.z46(q_10[18]),.z47(q_10[17]),.z48(q_10[16]),.z49(q_10[15]),.z50(q_10[14]),.z51(q_10[13]),.z52(q_10[12]),.z53(q_10[11]),.z54(q_10[10]),.z55(q_10[9]),.z56(q_10[8]),.z57(q_10[7]),.z58(q_10[6]),.z59(q_10[5]),.z60(q_10[4]),.z61(q_10[3]),.z62(q_10[2]),.z63(q_10[1]));

q_11 label11 ( .x0(X[64]),
.z00(q_11[64]),.z01(q_11[63]),.z02(q_11[62]),.z03(q_11[61]),.z04(q_11[60]),.z05(q_11[59]),.z06(q_11[58]),.z07(q_11[57]),.z08(q_11[56]),.z09(q_11[55]),.z10(q_11[54]),.z11(q_11[53]),.z12(q_11[52]),.z13(q_11[51]),.z14(q_11[50]),.z15(q_11[49]),.z16(q_11[48]),.z17(q_11[47]),.z18(q_11[46]),.z19(q_11[45]),.z20(q_11[44]),.z21(q_11[43]),.z22(q_11[42]),.z23(q_11[41]),.z24(q_11[40]),.z25(q_11[39]),.z26(q_11[38]),.z27(q_11[37]),.z28(q_11[36]),.z29(q_11[35]),.z30(q_11[34]),.z31(q_11[33]),.z32(q_11[32]),.z33(q_11[31]),.z34(q_11[30]),.z35(q_11[29]),.z36(q_11[28]),.z37(q_11[27]),.z38(q_11[26]),.z39(q_11[25]),.z40(q_11[24]),.z41(q_11[23]),.z42(q_11[22]),.z43(q_11[21]),.z44(q_11[20]),.z45(q_11[19]),.z46(q_11[18]),.z47(q_11[17]),.z48(q_11[16]),.z49(q_11[15]),.z50(q_11[14]),.z51(q_11[13]),.z52(q_11[12]),.z53(q_11[11]),.z54(q_11[10]),.z55(q_11[9]),.z56(q_11[8]),.z57(q_11[7]),.z58(q_11[6]),.z59(q_11[5]),.z60(q_11[4]),.z61(q_11[3]),.z62(q_11[2]),.z63(q_11[1]));


assign sum_res = X[3:1] + q_1[3:1] + q_2[3:1] + q_3[3:1]+ q_4[3:1]+ q_5[3:1] + q_6[3:1] + q_7[3:1] + q_8[3:1]+ q_9[3:1]+ q_10[3:1] + q_11[3:1];

quot_res  label12 (.x0(sum_res[6]),.x1(sum_res[5]),.x2(sum_res[4]),.x3(sum_res[3]),.x4(sum_res[2]),.x5(sum_res[1]),
                  .z0(sum[7]),.z1(sum[6]),.z2(sum[5]),.z3(sum[4]),.z4(sum[3]),.z5(sum[2]),.z6(sum[1]));

assign r_1 = q_1[9:4] + q_2[9:4] + q_3[9:4]+ q_4[9:4] + q_5[9:4] + q_6[9:4] + q_7[9:4] + q_8[9:4]+ q_9[9:4] + q_10[9:4] + q_11[9:4];

assign r_2 = r_1[10:7] + q_1[10] + q_2[15:10] + q_3[15:10] + q_4[15:10] + q_5[15:10] + q_6[15:10] + q_7[15:10] + q_8[15:10] + q_9[15:10] + q_10[15:10] + q_11[15:10];

assign r_3 = r_2[9:7] + q_2[16] + q_3[21:16] + q_4[21:16] + q_5[21:16] + q_6[21:16] + q_7[21:16] + q_8[21:16] + q_9[21:16] + q_10[21:16] + q_11[21:16];

assign r_4 = r_3[9:7] + q_3[22] + q_4[27:22] + q_5[27:22] + q_6[27:22] + q_7[27:22] + q_8[27:22] + q_9[27:22] + q_10[27:22] + q_11[27:22];

assign r_5 = r_4[9:7] + q_4[28] + q_5[33:28] + q_6[33:28] + q_7[33:28] + q_8[33:28] + q_9[33:28] + q_10[33:28] + q_11[33:28];

assign r_6 = r_5[9:7] + q_5[34] + q_6[39:34] + q_7[39:34] + q_8[39:34] + q_9[39:34] + q_10[39:34] + q_11[39:34];

assign r_7 = r_6[9:7] + q_6[40] + q_7[45:40] + q_8[45:40] + q_9[45:40] + q_10[45:40] + q_11[45:40];

assign r_8 = r_7[8:7] + q_7[46] + q_8[51:46] + q_9[51:46] + q_10[51:46] + q_11[51:46];

assign r_9 = r_8[8:7] + q_8[52] + q_9[57:52] + q_10[57:52] + q_11[57:52];

assign r_10 = r_9[8:7] + q_9[58] + q_10[63:58] + q_11[63:58];

assign r_11 = r_10[7] + q_10[64] + q_11[64];


assign Q = {r_11, r_10[6:1], r_9[6:1], r_8[6:1], r_7[6:1], r_6[6:1], r_5[6:1], r_4[6:1], r_3[6:1], r_2[6:1], r_1[6:1]} + sum[7:4];

assign R = sum[3:1]; 

endmodule