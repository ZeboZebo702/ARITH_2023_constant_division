// Benchmark "q_4" written by ABC on Tue Jul 04 13:16:23 2023

module q_4 ( 
    x0, x1, x2, x3, x4, x5,
    z0, z1, z2, z3, z4  );
  input  x0, x1, x2, x3, x4, x5;
  output z0, z1, z2, z3, z4;
  assign z0 = (x4 & ((x0 & x1 & ~x2 & x3) | (~x0 & ~x1 & x2 & ~x3))) | (~x4 & (x0 ? (x1 ? (x2 & ~x3) : (~x2 ^ x3)) : (x1 ? (~x2 & x3) : (x2 & ~x3)))) | (x4 & (~x2 ^ x5) & (x0 ? (~x1 & ~x3) : (x1 & x3)));
  assign z1 = (~x2 & ((x1 & (x0 ? (x3 ^ x4) : ~x3)) | (~x0 & ~x1 & x3))) | (x2 & ((x0 & (x1 ? (x3 & x4) : (~x3 & ~x4))) | (x3 & ~x4 & ~x0 & x1))) | (x4 & (x0 ? (~x1 & (x2 ? (~x3 & ~x5) : (x3 & x5))) : (x1 & x2 & (x3 ^ x5))));
  assign z2 = ((x4 ^ x5) & ((~x0 & x1 & x2) | (x0 & ~x1 & ~x2) | (x2 & ~x3 & x0 & ~x1))) | (~x0 & ~x1 & x4) | (x0 & x1 & ~x4) | (~x0 & x1 & ~x2 & ~x3 & x4) | (x3 & ((x0 & ~x1 & x2 & ~x4 & x5) | (~x0 & x1 & ~x2 & x4 & ~x5)));
  assign z3 = (~x5 & (x0 ? (~x1 & ~x2) : (x1 & x2))) | (x5 & (~x0 ^ x1)) | (~x3 & ((~x0 & x1 & ~x2 & x5) | (x0 & ~x1 & x2 & ~x5))) | (x3 & ((x0 & ~x1 & x2 & (~x4 ^ x5)) | (~x0 & x1 & ~x2 & ~x4 & x5)));
  assign z4 = (~x0 & (x1 ? (~x2 & ~x3) : (x2 & x3))) | (x0 & (x1 ? (x2 & x3) : (x2 ^ x3))) | (x0 & x2 & (x1 ? (~x3 & x4) : (x3 & ~x4))) | (~x0 & x1 & ~x2 & x3 & ~x4) | (~x2 & x4 & ((~x3 & x5 & x0 & ~x1) | (~x0 & x1 & x3 & ~x5)));
endmodule


