module div_48_113(X, Q, R );

input  [48:1] X;
output [42:1] Q;  
output [7:1] R;  

wire [42:1] Q_temp;
wire [10:1] r_1;
wire [10:1] r_2;
wire [9:1] r_3;
wire [9:1] r_4;
wire [8:1] r_5;
wire [7:1] r_6;


wire [10:1] sum_res;
wire [10:1] sum;

wire [15:1] q_1;
wire [22:1] q_2;
wire [29:1] q_3;
wire [36:1] q_4;
wire [43:1] q_5;
wire [49:1] q_6;


q_1 label1 ( .x0(X[14]),.x1(X[13]),.x2(X[12]),.x3(X[11]),.x4(X[10]),.x5(X[9]),.x6(X[8]),
.z00(q_1[15]),.z01(q_1[14]),.z02(q_1[13]),.z03(q_1[12]),.z04(q_1[11]),.z05(q_1[10]),.z06(q_1[9]),.z07(q_1[8]),.z08(q_1[7]),.z09(q_1[6]),.z10(q_1[5]),.z11(q_1[4]),.z12(q_1[3]),.z13(q_1[2]),.z14(q_1[1]));

q_2 label2 ( .x0(X[21]),.x1(X[20]),.x2(X[19]),.x3(X[18]),.x4(X[17]),.x5(X[16]),.x6(X[15]),
.z00(q_2[22]),.z01(q_2[21]),.z02(q_2[20]),.z03(q_2[19]),.z04(q_2[18]),.z05(q_2[17]),.z06(q_2[16]),.z07(q_2[15]),.z08(q_2[14]),.z09(q_2[13]),.z10(q_2[12]),.z11(q_2[11]),.z12(q_2[10]),.z13(q_2[9]),.z14(q_2[8]),.z15(q_2[7]),.z16(q_2[6]),.z17(q_2[5]),.z18(q_2[4]),.z19(q_2[3]),.z20(q_2[2]),.z21(q_2[1]));

q_3 label3 ( .x0(X[28]),.x1(X[27]),.x2(X[26]),.x3(X[25]),.x4(X[24]),.x5(X[23]),.x6(X[22]),
.z00(q_3[29]),.z01(q_3[28]),.z02(q_3[27]),.z03(q_3[26]),.z04(q_3[25]),.z05(q_3[24]),.z06(q_3[23]),.z07(q_3[22]),.z08(q_3[21]),.z09(q_3[20]),.z10(q_3[19]),.z11(q_3[18]),.z12(q_3[17]),.z13(q_3[16]),.z14(q_3[15]),.z15(q_3[14]),.z16(q_3[13]),.z17(q_3[12]),.z18(q_3[11]),.z19(q_3[10]),.z20(q_3[9]),.z21(q_3[8]),.z22(q_3[7]),.z23(q_3[6]),.z24(q_3[5]),.z25(q_3[4]),.z26(q_3[3]),.z27(q_3[2]),.z28(q_3[1]));

q_4 label4 ( .x0(X[35]),.x1(X[34]),.x2(X[33]),.x3(X[32]),.x4(X[31]),.x5(X[30]),.x6(X[29]),
.z00(q_4[36]),.z01(q_4[35]),.z02(q_4[34]),.z03(q_4[33]),.z04(q_4[32]),.z05(q_4[31]),.z06(q_4[30]),.z07(q_4[29]),.z08(q_4[28]),.z09(q_4[27]),.z10(q_4[26]),.z11(q_4[25]),.z12(q_4[24]),.z13(q_4[23]),.z14(q_4[22]),.z15(q_4[21]),.z16(q_4[20]),.z17(q_4[19]),.z18(q_4[18]),.z19(q_4[17]),.z20(q_4[16]),.z21(q_4[15]),.z22(q_4[14]),.z23(q_4[13]),.z24(q_4[12]),.z25(q_4[11]),.z26(q_4[10]),.z27(q_4[9]),.z28(q_4[8]),.z29(q_4[7]),.z30(q_4[6]),.z31(q_4[5]),.z32(q_4[4]),.z33(q_4[3]),.z34(q_4[2]),.z35(q_4[1]));

q_5 label5 ( .x0(X[42]),.x1(X[41]),.x2(X[40]),.x3(X[39]),.x4(X[38]),.x5(X[37]),.x6(X[36]),
.z00(q_5[43]),.z01(q_5[42]),.z02(q_5[41]),.z03(q_5[40]),.z04(q_5[39]),.z05(q_5[38]),.z06(q_5[37]),.z07(q_5[36]),.z08(q_5[35]),.z09(q_5[34]),.z10(q_5[33]),.z11(q_5[32]),.z12(q_5[31]),.z13(q_5[30]),.z14(q_5[29]),.z15(q_5[28]),.z16(q_5[27]),.z17(q_5[26]),.z18(q_5[25]),.z19(q_5[24]),.z20(q_5[23]),.z21(q_5[22]),.z22(q_5[21]),.z23(q_5[20]),.z24(q_5[19]),.z25(q_5[18]),.z26(q_5[17]),.z27(q_5[16]),.z28(q_5[15]),.z29(q_5[14]),.z30(q_5[13]),.z31(q_5[12]),.z32(q_5[11]),.z33(q_5[10]),.z34(q_5[9]),.z35(q_5[8]),.z36(q_5[7]),.z37(q_5[6]),.z38(q_5[5]),.z39(q_5[4]),.z40(q_5[3]),.z41(q_5[2]),.z42(q_5[1]));

q_6 label6 ( .x0(X[48]),.x1(X[47]),.x2(X[46]),.x3(X[45]),.x4(X[44]),.x5(X[43]),
.z00(q_6[49]),.z01(q_6[48]),.z02(q_6[47]),.z03(q_6[46]),.z04(q_6[45]),.z05(q_6[44]),.z06(q_6[43]),.z07(q_6[42]),.z08(q_6[41]),.z09(q_6[40]),.z10(q_6[39]),.z11(q_6[38]),.z12(q_6[37]),.z13(q_6[36]),.z14(q_6[35]),.z15(q_6[34]),.z16(q_6[33]),.z17(q_6[32]),.z18(q_6[31]),.z19(q_6[30]),.z20(q_6[29]),.z21(q_6[28]),.z22(q_6[27]),.z23(q_6[26]),.z24(q_6[25]),.z25(q_6[24]),.z26(q_6[23]),.z27(q_6[22]),.z28(q_6[21]),.z29(q_6[20]),.z30(q_6[19]),.z31(q_6[18]),.z32(q_6[17]),.z33(q_6[16]),.z34(q_6[15]),.z35(q_6[14]),.z36(q_6[13]),.z37(q_6[12]),.z38(q_6[11]),.z39(q_6[10]),.z40(q_6[9]),.z41(q_6[8]),.z42(q_6[7]),.z43(q_6[6]),.z44(q_6[5]),.z45(q_6[4]),.z46(q_6[3]),.z47(q_6[2]),.z48(q_6[1]));


assign sum_res = X[7:1] + q_1[7:1] + q_2[7:1] + q_3[7:1] + q_4[7:1] + q_5[7:1] + q_6[7:1];

quot_res  label9 (.x0(sum_res[10]),.x1(sum_res[9]),.x2(sum_res[8]),.x3(sum_res[7]),.x4(sum_res[6]),.x5(sum_res[5]),.x6(sum_res[4]),
		  .x7(sum_res[3]),.x8(sum_res[2]),.x9(sum_res[1]),
                  .z0(sum[10]),.z1(sum[9]),.z2(sum[8]),.z3(sum[7]),.z4(sum[6]),.z5(sum[5]),
		  .z6(sum[4]),.z7(sum[3]),.z8(sum[2]),.z9(sum[1]));

assign r_1 = q_1[14:8] + q_2[14:8] + q_3[14:8] + q_4[14:8] + q_5[14:8] + q_6[14:8];

assign r_2 = q_1[15] + r_1[10:8] + q_2[21:15] + q_3[21:15] + q_4[21:15] + q_5[21:15] + q_6[21:15];

assign r_3 = r_2[10:8] + q_2[22] + q_3[28:22] + q_4[28:22] + q_5[28:22] + q_6[28:22];

assign r_4 = r_3[9:8] + q_3[29] + q_4[35:29] + q_5[35:29] + q_6[35:29];

assign r_5 = r_4[9:8] + q_4[36] + q_5[42:36] + q_6[42:36];

assign r_6 = r_5[8] + q_5[43] + q_6[49:43];


assign Q_temp = {r_6[7:1], r_5[7:1], r_4[7:1], r_3[7:1], r_2[7:1], r_1[7:1]};

assign Q = Q_temp + sum[10:8];

assign R = sum[7:1]; 

endmodule