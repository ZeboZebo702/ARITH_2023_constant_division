module div_32_3(X, Q, R );

input  [32:1] X;
output [31:1] Q;  
output [2:1] R;  

//wire [28:1] Q_temp;

wire [8:1] r_1;
wire [8:1] r_2;
wire [7:1] r_3;
wire [7:1] r_4;
wire [6:1] r_5;

wire [4:1] sum_res;
wire [5:1] sum;

wire [7:1] q_1;
wire [13:1] q_2;
wire [19:1] q_3;
wire [25:1] q_4;
wire [31:1] q_5;


q_1 label1 ( .x0(X[8]),.x1(X[7]),.x2(X[6]),.x3(X[5]),.x4(X[4]),.x5(X[3]),
.z0(q_1[7]),.z1(q_1[6]),.z2(q_1[5]),.z3(q_1[4]),.z4(q_1[3]),.z5(q_1[2]),.z6(q_1[1]));

q_2 label2 ( .x0(X[14]),.x1(X[13]),.x2(X[12]),.x3(X[11]),.x4(X[10]),.x5(X[9]),
.z00(q_2[13]),.z01(q_2[12]),.z02(q_2[11]),.z03(q_2[10]),.z04(q_2[9]),.z05(q_2[8]),.z06(q_2[7]),.z07(q_2[6]),.z08(q_2[5]),.z09(q_2[4]),.z10(q_2[3]),.z11(q_2[2]),.z12(q_2[1]));

q_3 label3 ( .x0(X[20]),.x1(X[19]),.x2(X[18]),.x3(X[17]),.x4(X[16]),.x5(X[15]),
.z00(q_3[19]),.z01(q_3[18]),.z02(q_3[17]),.z03(q_3[16]),.z04(q_3[15]),.z05(q_3[14]),.z06(q_3[13]),.z07(q_3[12]),.z08(q_3[11]),.z09(q_3[10]),.z10(q_3[9]),.z11(q_3[8]),.z12(q_3[7]),.z13(q_3[6]),.z14(q_3[5]),.z15(q_3[4]),.z16(q_3[3]),.z17(q_3[2]),.z18(q_3[1]));

q_4 label4 ( .x0(X[26]),.x1(X[25]),.x2(X[24]),.x3(X[23]),.x4(X[22]),.x5(X[21]),
.z00(q_4[25]),.z01(q_4[24]),.z02(q_4[23]),.z03(q_4[22]),.z04(q_4[21]),.z05(q_4[20]),.z06(q_4[19]),.z07(q_4[18]),.z08(q_4[17]),.z09(q_4[16]),.z10(q_4[15]),.z11(q_4[14]),.z12(q_4[13]),.z13(q_4[12]),.z14(q_4[11]),.z15(q_4[10]),.z16(q_4[9]),.z17(q_4[8]),.z18(q_4[7]),.z19(q_4[6]),.z20(q_4[5]),.z21(q_4[4]),.z22(q_4[3]),.z23(q_4[2]),.z24(q_4[1]));

q_5 label5 ( .x0(X[32]),.x1(X[31]),.x2(X[30]),.x3(X[29]),.x4(X[28]),.x5(X[27]),
.z00(q_5[31]),.z01(q_5[30]),.z02(q_5[29]),.z03(q_5[28]),.z04(q_5[27]),.z05(q_5[26]),.z06(q_5[25]),.z07(q_5[24]),.z08(q_5[23]),.z09(q_5[22]),.z10(q_5[21]),.z11(q_5[20]),.z12(q_5[19]),.z13(q_5[18]),.z14(q_5[17]),.z15(q_5[16]),.z16(q_5[15]),.z17(q_5[14]),.z18(q_5[13]),.z19(q_5[12]),.z20(q_5[11]),.z21(q_5[10]),.z22(q_5[9]),.z23(q_5[8]),.z24(q_5[7]),.z25(q_5[6]),.z26(q_5[5]),.z27(q_5[4]),.z28(q_5[3]),.z29(q_5[2]),.z30(q_5[1]));


assign sum_res = X[2:1] + q_1[2:1] + q_2[2:1] + q_3[2:1] + q_4[2:1] + q_5[2:1];

quot_res  label10 (.x0(sum_res[4]),.x1(sum_res[3]),.x2(sum_res[2]),.x3(sum_res[1]),
                  .z0(sum[5]),.z1(sum[4]),.z2(sum[3]),.z3(sum[2]),.z4(sum[1]));


assign r_1 = q_1[6:1] + q_2[6:1] + q_3[6:1] + q_4[6:1] + q_5[6:1];

assign r_2 = r_1[8:7] + q_1[7] + q_2[12:7] + q_3[12:7] + q_4[12:7] + q_5[12:7];

assign r_3 = r_2[8:7] + q_2[13] + q_3[18:13] + q_4[18:13] + q_5[18:13];

assign r_4 = r_3[7] + q_3[19] + q_4[24:19] + q_5[24:19];

assign r_5 = r_4[7] + q_4[25] + q_5[30:25];

assign Q = {q_5[31], r_5[6:1], r_4[6:1], r_3[6:1], r_2[6:1], r_1[6:1]} + sum[5:3];


//assign Q = Q_temp;

assign R = sum[2:1]; 

endmodule