module div_38_47(X, Q, R );

input  [36:0] X;
output [31:1] Q;  
output [6:1] R;  

wire [31:1] Q_temp;
wire [9:1] r_1;
wire [8:1] r_2;
wire [8:1] r_3;
wire [7:1] r_4;
wire [6:1] r_5;

wire [9:1] sum_res;
wire [9:1] sum;

wire [13:1] q_1;
wire [19:1] q_2;
wire [25:1] q_3;
wire [31:1] q_4;
wire [37:1] q_5;

q_1 label1 ( .x0(X[12]),.x1(X[11]),.x2(X[10]),.x3(X[9]),.x4(X[8]),.x5(X[7]),
.z00(q_1[13]),.z01(q_1[12]),.z02(q_1[11]),.z03(q_1[10]),.z04(q_1[9]),.z05(q_1[8]),.z06(q_1[7]),.z07(q_1[6]),.z08(q_1[5]),.z09(q_1[4]),.z10(q_1[3]),.z11(q_1[2]),.z12(q_1[1]));

q_2 label2 ( .x0(X[18]),.x1(X[17]),.x2(X[16]),.x3(X[15]),.x4(X[14]),.x5(X[13]),
.z00(q_2[19]),.z01(q_2[18]),.z02(q_2[17]),.z03(q_2[16]),.z04(q_2[15]),.z05(q_2[14]),.z06(q_2[13]),.z07(q_2[12]),.z08(q_2[11]),.z09(q_2[10]),.z10(q_2[9]),.z11(q_2[8]),.z12(q_2[7]),.z13(q_2[6]),.z14(q_2[5]),.z15(q_2[4]),.z16(q_2[3]),.z17(q_2[2]),.z18(q_2[1]));

q_3 label3 ( .x0(X[24]),.x1(X[23]),.x2(X[22]),.x3(X[21]),.x4(X[20]),.x5(X[19]),
.z00(q_3[25]),.z01(q_3[24]),.z02(q_3[23]),.z03(q_3[22]),.z04(q_3[21]),.z05(q_3[20]),.z06(q_3[19]),.z07(q_3[18]),.z08(q_3[17]),.z09(q_3[16]),.z10(q_3[15]),.z11(q_3[14]),.z12(q_3[13]),.z13(q_3[12]),.z14(q_3[11]),.z15(q_3[10]),.z16(q_3[9]),.z17(q_3[8]),.z18(q_3[7]),.z19(q_3[6]),.z20(q_3[5]),.z21(q_3[4]),.z22(q_3[3]),.z23(q_3[2]),.z24(q_3[1]));

q_4 label4 ( .x0(X[30]),.x1(X[29]),.x2(X[28]),.x3(X[27]),.x4(X[26]),.x5(X[25]),
.z00(q_4[31]),.z01(q_4[30]),.z02(q_4[29]),.z03(q_4[28]),.z04(q_4[27]),.z05(q_4[26]),.z06(q_4[25]),.z07(q_4[24]),.z08(q_4[23]),.z09(q_4[22]),.z10(q_4[21]),.z11(q_4[20]),.z12(q_4[19]),.z13(q_4[18]),.z14(q_4[17]),.z15(q_4[16]),.z16(q_4[15]),.z17(q_4[14]),.z18(q_4[13]),.z19(q_4[12]),.z20(q_4[11]),.z21(q_4[10]),.z22(q_4[9]),.z23(q_4[8]),.z24(q_4[7]),.z25(q_4[6]),.z26(q_4[5]),.z27(q_4[4]),.z28(q_4[3]),.z29(q_4[2]),.z30(q_4[1]));

q_5 label5 ( .x0(X[36]),.x1(X[35]),.x2(X[34]),.x3(X[33]),.x4(X[32]),.x5(X[31]),
.z00(q_5[37]),.z01(q_5[36]),.z02(q_5[35]),.z03(q_5[34]),.z04(q_5[33]),.z05(q_5[32]),.z06(q_5[31]),.z07(q_5[30]),.z08(q_5[29]),.z09(q_5[28]),.z10(q_5[27]),.z11(q_5[26]),.z12(q_5[25]),.z13(q_5[24]),.z14(q_5[23]),.z15(q_5[22]),.z16(q_5[21]),.z17(q_5[20]),.z18(q_5[19]),.z19(q_5[18]),.z20(q_5[17]),.z21(q_5[16]),.z22(q_5[15]),.z23(q_5[14]),.z24(q_5[13]),.z25(q_5[12]),.z26(q_5[11]),.z27(q_5[10]),.z28(q_5[9]),.z29(q_5[8]),.z30(q_5[7]),.z31(q_5[6]),.z32(q_5[5]),.z33(q_5[4]),.z34(q_5[3]),.z35(q_5[2]),.z36(q_5[1]));

assign sum_res = X[6:1] + q_1[6:1] + q_2[6:1] + q_3[6:1] + q_4[6:1] + q_5[6:1];

quot_res  label10 (.x0(sum_res[9]),.x1(sum_res[8]),.x2(sum_res[7]),.x3(sum_res[6]),.x4(sum_res[5]),
		  .x5(sum_res[4]),.x6(sum_res[3]),.x7(sum_res[2]),.x8(sum_res[1]),
                  .z0(sum[9]),.z1(sum[8]),.z2(sum[7]),.z3(sum[6]),.z4(sum[5]),
		  .z5(sum[4]),.z6(sum[3]),.z7(sum[2]),.z8(sum[1]));


assign r_1 = q_1[12:7] + q_2[12:7] + q_3[12:7] + q_4[12:7] + q_5[12:7];

assign r_2 = r_1[9:7] + q_1[13] + q_2[18:13] + q_3[18:13] + q_4[18:13] + q_5[18:13];

assign r_3 = r_2[8:7] + q_2[19] + q_3[24:19] + q_4[24:19] + q_5[24:19];

assign r_4 = r_3[8:7] + q_3[25] + q_4[30:25] + q_5[30:25];

assign r_5 = r_4[7] + q_4[31] + q_5[36:31];

assign Q_temp = {r_5[6:1], r_4[6:1], r_3[6:1], r_2[6:1], r_1[6:1]};


assign Q = Q_temp + sum[9:7];

assign R = sum[6:1]; 

endmodule