// Benchmark "quot_res" written by ABC on Fri Feb 24 17:34:06 2023

module quot_res ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10;
  wire n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n36, n37, n38,
    n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n50, n51, n52, n53,
    n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
    n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n81, n82,
    n83, n84, n85, n86, n87, n89, n90, n91, n92, n93, n94, n95, n96, n97,
    n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
    n110, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n152, n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n257, n258,
    n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
    n283, n284, n285, n286, n287, n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302, n303;
  assign z00 = n24 | ~n25 | n27 | n31 | n33;
  assign n24 = x04 & ((x00 & (~x01 | ~x02 | (~x03 & ~x05))) | (~x00 & x01 & x02 & x03 & x05));
  assign n25 = (x00 | ~x01 | ~x02 | ~x03 | ~n26) & (~x00 | x04 | (x01 & x02 & x03));
  assign n26 = x07 & ~x06 & x04 & ~x05;
  assign n27 = n30 & n28 & n29;
  assign n28 = x04 & ~x03 & x02 & x00 & x01;
  assign n29 = x05 & x06;
  assign n30 = ~x09 & ~x07 & ~x08;
  assign n31 = ~n32 & x04 & x01 & x02;
  assign n32 = (~x00 | x03 | ~x05 | x06) & (x00 | ~x03 | x05 | ~x06);
  assign n33 = n34 & x08 & ~x06 & ~x07;
  assign n34 = ~x05 & x04 & x03 & ~x00 & x01 & x02;
  assign z01 = n43 | ~n44 | (n41 & (~n42 | (~x07 & ~n36)));
  assign n36 = (~x00 | n37) & (x00 | ~n38 | ~n39 | ~n40);
  assign n37 = (~x01 | x03 | ~x04 | ~x06 | x08 | x09) & (x01 | ~x03 | x04 | x06 | ~x08 | ~x09);
  assign n38 = ~x01 & x03;
  assign n39 = x04 & ~x06;
  assign n40 = ~x08 & x09;
  assign n41 = x02 & x05;
  assign n42 = (~x00 | ((x01 | ~x03 | x04 | ~x06) & (~x01 | x03 | ~x04 | x06))) & (x00 | x01 | ~x03 | ~x04 | ~x06);
  assign n43 = x00 & ((x01 & (~x02 | (~x03 & ~x04))) | (x03 & x04 & ~x01 & x02));
  assign n44 = ~n47 & n45 & (x06 | ~n38 | ~n41 | ~n46);
  assign n45 = ~x01 | ((x03 | (x00 & (~x02 | ~x04 | x05))) & (x00 | (x02 & x04)));
  assign n46 = x07 & (x00 ^ x04);
  assign n47 = n48 & (x01 ? (~x05 & ~x08) : (x05 & x08));
  assign n48 = ~x07 & ~x06 & x04 & ~x00 & x02 & x03;
  assign z02 = ~n68 | ~n65 | ~n61 | n50 | n56;
  assign n50 = n55 & ((n53 & n54) | (n51 & ~n52));
  assign n51 = ~x00 & x04;
  assign n52 = (x01 | x02 | ~x05 | ~x06 | ~x08) & (~x01 | x05 | (x02 ? (x06 | x08) : (~x06 | ~x08)));
  assign n53 = x02 & x00 & ~x01;
  assign n54 = ~x04 & x05 & ~x06 & ~x08;
  assign n55 = x03 & ~x07;
  assign n56 = x05 & ~x07 & ((~n57 & n58) | (n59 & n60));
  assign n57 = x00 ? (x04 | ~x08) : (~x04 | x08);
  assign n58 = ~x01 & x03 & (x02 ? (~x06 & ~x09) : (x06 & x09));
  assign n59 = ~x03 & x02 & x00 & x01;
  assign n60 = ~x09 & ~x08 & x04 & x06;
  assign n61 = ~n64 & (~x00 | ~x02 | ~n62 | (x01 & ~n63));
  assign n62 = ~x03 & x04;
  assign n63 = x05 & ~x06;
  assign n64 = ~x05 & x04 & ~x03 & x02 & x00 & x01;
  assign n65 = ~x03 | n66 | ((x02 | ((~x05 | ~n67) & (~x01 | (~x05 & ~n67)))) & (x01 | ~x02 | x05));
  assign n66 = ~x00 ^ x04;
  assign n67 = x06 & x07;
  assign n68 = n70 & (~x10 | ~n69 | ~n71 | ~n72);
  assign n69 = ~x02 & x03;
  assign n70 = (~x02 | ((x00 | (x03 & x04)) & (x03 | x04))) & (~x03 | ~x04 | ~x00 | x02);
  assign n71 = (x01 ? (~x05 & x09) : (x05 & ~x09)) & (x00 ? (~x04 & x08) : (x04 & ~x08));
  assign n72 = x06 & ~x07;
  assign z03 = ~n79 | (x07 ? (~x03 & ~n84) : (~n74 | ~n85));
  assign n74 = ~n75 & (~n51 | n78);
  assign n75 = x00 & (x01 ? (n69 & n77) : ~n76);
  assign n76 = (x02 | ((x03 | ~x04 | x05 | x06 | ~x08) & (~x03 | x04 | ~x05 | ~x06 | x08))) & (~x05 | x06 | x08 | ~x02 | ~x03 | x04);
  assign n77 = ~x08 & x06 & ~x04 & ~x05;
  assign n78 = (x03 | ~x08 | ((~x01 | (x02 ? (x05 | ~x06) : (~x05 | x06))) & (x01 | ~x02 | ~x05 | ~x06))) & (~x01 | ~x02 | ~x03 | x05 | x06 | x08);
  assign n79 = ~n81 & n82 & n83 & (x02 | n80);
  assign n80 = (((~x01 | (x03 ? (x05 | x06) : (~x05 | ~x06))) & (x01 | ~x03 | ~x05 | x06)) | (~x00 ^ x04)) & (~x00 | x01 | x03 | ~x04 | x05 | ~x06);
  assign n81 = n71 & n72 & (x02 ? (~x03 & x10) : (x03 & ~x10));
  assign n82 = x00 ? (x03 | ~x04 | (x02 ? (x01 & ~n63) : ~x01)) : (~x03 | x04);
  assign n83 = (((x01 | ~x03 | x05) & (~x01 | ~x02 | x03 | ~x05)) | (~x00 ^ x04)) & (~x00 | x03 | ~x04 | (x01 ? (~x02 | x05) : (x02 | ~x05)));
  assign n84 = ((~x00 ^ x04) | ((~x01 | (x02 ? (x05 | ~x06) : (~x05 | x06))) & (x01 | ~x02 | ~x05 | ~x06))) & (~x04 | x05 | x06 | ~x00 | x01 | x02);
  assign n85 = (~n59 | ~n87) & (n57 | n86);
  assign n86 = x01 ? (x02 | ((x03 | ~x05 | x06 | ~x09) & (~x03 | x05 | ~x06 | x09))) : (~x02 | ~x05 | (x03 ? (x06 | x09) : (~x06 | ~x09)));
  assign n87 = ~x09 & ~x08 & x06 & x04 & x05;
  assign z04 = n101 | ~n104 | (~x07 & (~n89 | n94 | n98));
  assign n89 = (x05 | n90) & (x04 | ~x05 | n93);
  assign n90 = (x06 | n91) & (~x01 | x04 | ~x06 | n92);
  assign n91 = (~x00 | x01 | x02 | ((x04 | ~x08) & (x03 | ~x04 | x08))) & (x00 | ~x01 | ~x02 | ~x03 | ~x04 | x08);
  assign n92 = x00 ? (x08 | (~x02 ^ x03)) : (~x02 | ~x08);
  assign n93 = ((x01 ? (x02 | x06) : (~x02 | ~x06)) | (x00 ? (x03 | x08) : ~x08)) & (~x00 | x01 | ~x03 | x08 | (~x02 ^ x06));
  assign n94 = x06 & ((~n95 & ~n96) | (~x08 & n41 & ~n97));
  assign n95 = ~x02 ^ x03;
  assign n96 = (~x00 | ~x08 | ((~x05 | ~x09 | x01 | ~x04) & (x05 | x09 | ~x01 | x04))) & (x00 | ~x01 | ~x04 | x05 | x08 | x09);
  assign n97 = (x00 | x01 | x04 | ~x09) & (~x00 | ~x01 | x03 | ~x04 | x09);
  assign n98 = n63 & (n100 | (~n99 & (x01 ? (~x02 & ~x03) : (x02 & x03))));
  assign n99 = (~x00 | ~x08 | (~x04 ^ ~x09)) & (x00 | ~x04 | x08 | x09);
  assign n100 = ~x00 & x01 & ~x02 & ~x04 & ~x08 & x09;
  assign n101 = x07 & (n102 | (x00 & x04 & ~n103));
  assign n102 = ~x04 & ((~x00 & ((x01 & (x02 ? (~x05 & x06) : (x05 & ~x06))) | (~x01 & x02 & x05 & x06))) | (x00 & ~x01 & ~x02 & ~x05 & ~x06));
  assign n103 = (~x06 | (~x01 ^ x05) | (~x02 ^ x03)) & (~x05 | x06 | (x01 ? (x02 | x03) : (~x02 | ~x03)));
  assign n104 = ~n106 & ~n107 & ~n109 & (x06 ? n105 : n110);
  assign n105 = (x02 | ((~x00 | ((~x04 | ~x05 | ~x01 | x03) & (x01 | x04 | x05))) & (x00 | ~x01 | x04 | ~x05))) & (~x00 | x01 | ~x02 | ~x03 | ~x04 | ~x05);
  assign n106 = ~x02 & (x00 ? ((x01 & (x03 ? (x04 & x05) : (~x04 & ~x05))) | (~x01 & ~x03 & ~x04 & x05)) : (x04 & ((~x03 & ~x05) | (~x01 & (~x03 | ~x05)))));
  assign n107 = n72 & ~n108 & (x01 ? (~x05 & x09) : (x05 & ~x09));
  assign n108 = x02 ? ((x03 | ((~x00 | ~x08 | (~x04 ^ ~x10)) & (x08 | x10 | x00 | ~x04))) & (x08 | ~x10 | x00 | x04)) : (~x03 | ((~x00 | ~x08 | (~x04 ^ ~x10)) & (x08 | x10 | x00 | ~x04)));
  assign n109 = x02 & ((~x00 & (x01 ? (~x04 & x05) : (x04 & ~x05))) | (x00 & ~x01 & ~x04 & ~x05));
  assign n110 = (x00 & x04 & (~x01 | ~x05)) | (~x00 & (~x04 | (x01 & x05))) | (x01 & x05 & (x03 | ~x04)) | (x02 & x03) | (~x02 & ~x03) | (~x01 & ~x05);
  assign z05 = n112 | ~n124 | ~n137 | ~n145 | (~x03 & ~n123);
  assign n112 = n72 & (~n118 | (x02 & (n116 | (~x03 & ~n113))));
  assign n113 = (x01 | x09 | n114) & (~x00 | ~x01 | ~x04 | ~n115);
  assign n114 = (~x00 | ~x08 | ((x05 | ~x10) & (~x04 | ~x05 | x10))) & (x08 | ~x10 | x00 | x05);
  assign n115 = ~x10 & ~x05 & x08 & x09;
  assign n116 = n117 & (x00 ? (~x04 & x08) : ~x08);
  assign n117 = ~x01 & x03 & ~x05 & ~x09 & x10;
  assign n118 = (~n121 | ~n122) & (n119 | n120);
  assign n119 = (~x01 | ~x09 | (~x05 ^ ~x10)) & (x01 | ~x05 | x09 | x10);
  assign n120 = x00 ? (~x08 | (x02 ? (x03 | x04) : ~x03)) : (x08 | (x02 ^ (~x03 | ~x04)));
  assign n121 = x08 & x00 & ~x01;
  assign n122 = x10 & ~x09 & ~x05 & ~x02 & x03 & x04;
  assign n123 = (x02 | ((x00 | x01 | ~x05) & (~x00 | ~x01 | x05 | ~x06))) & (~x01 | ((~x00 | x05 | x06 | (~x02 & ~x07)) & (x00 | ~x02 | ~x05 | ~x06 | ~x07))) & (x01 | ((x00 | ~x05 | x06) & (~x02 | x05 | ~x06 | ~x07)));
  assign n124 = n125 & ~n129 & (~n55 | (~n132 & ~n134));
  assign n125 = (~x00 | (x01 ? (~n126 | ~n128) : (~x05 | n127))) & (x00 | ~x01 | x05 | n127);
  assign n126 = x02 & ~x03;
  assign n127 = (x06 & (x02 | x03)) | (x02 & x03 & (x07 | x08)) | (~x07 & ~x08 & ~x02 & ~x06);
  assign n128 = x07 & ~x04 & x05 & x06;
  assign n129 = ~x07 & (x01 ? (x05 ? ~n130 : (~n95 & n131)) : (x05 ? (~n95 & n131) : ~n130));
  assign n130 = (x00 | ~x02 | ~x06 | ~x08) & (~x00 | x02 | x03 | x06 | x08);
  assign n131 = ~x08 & x00 & x06;
  assign n132 = ~x06 & ~n133 & (x01 ? (~x02 & ~x09) : (x02 & x09));
  assign n133 = (x00 | x04 | ~x05 | x08) & (~x00 | ~x04 | x05 | ~x08);
  assign n134 = n135 & ~n136 & (x02 ^ x09);
  assign n135 = ~x05 & x06;
  assign n136 = (~x04 | ~x08 | ~x00 | x01) & (x00 | ~x01 | x04 | x08);
  assign n137 = (n138 | ~n139) & (~n55 | (~n140 & n142));
  assign n138 = (~x02 | ((x01 | ((x05 | ~x06 | ~x09) & (~x03 | ~x05 | x06 | x09))) & (~x01 | x03 | x05 | ~x06 | x09))) & (~x01 | x02 | ((x05 | ((~x03 | ~x06 | x09) & (x06 | ~x09))) & (x03 | ~x05 | x06 | x09)));
  assign n139 = ~x07 & (x00 ^ ~x08);
  assign n140 = ~n141 & x04 & ~x08;
  assign n141 = (~x00 | x05 | (x01 ? (x02 | x06) : (~x02 | ~x06))) & (x00 | ~x01 | ~x02 | ~x05 | ~x06);
  assign n142 = x04 ? (~x05 | n143) : ((x05 | n143) & (~x08 | ~n144 | ~x05 | x06));
  assign n143 = (~x00 | x01 | x02 | x06 | x08) & (x00 | ~x01 | ~x08 | (x02 ^ ~x06));
  assign n144 = x02 & ~x00 & ~x01;
  assign n145 = ~x03 | (n147 & (n148 | ~n149) & (~n146 | ~n150));
  assign n146 = ~x02 & ~x00 & ~x01;
  assign n147 = (~x07 | ((x01 | ~x02 | x05 | ~x06) & (~x01 | ((x00 | ~x02 | ~x05 | ~x06) & (~x00 | x02 | (x05 ^ x06)))))) & (x00 | x01 | x02 | ~x05 | x06);
  assign n148 = (~x00 | x01 | ~x04 | x05) & (x00 | (x01 ? (x04 ^ x05) : (x04 | ~x05)));
  assign n149 = x07 & (x02 ^ x06);
  assign n150 = ~x07 & ~x04 & x05 & x06;
  assign z06 = n152 | n157 | ~n159 | n175 | (~x07 & ~n177);
  assign n152 = x04 & (n155 | (x02 & (n154 | (~x07 & ~n153))));
  assign n153 = (~x01 | x08 | ((x05 | ~x06 | ~x00 | x03) & (x00 | ~x03 | ~x05 | x06))) & (x00 | x01 | ~x03 | ~x08 | (x05 ^ x06));
  assign n154 = ~x00 & ~x01 & x03 & x07 & (~x05 ^ x06);
  assign n155 = ~n156 & x03 & ~x00 & ~x02;
  assign n156 = x01 ? (~x05 | x06 | (~x07 & ~x08)) : (x05 | ~x06);
  assign n157 = ~n158 & ~x04 & x00 & x03;
  assign n158 = ((x01 ? (x02 | ~x05) : (~x02 | x05)) | (x06 ? (x07 | x08) : ~x07)) & (x01 | ~x06 | (x02 ? (~x05 | ~x07) : (x05 | (~x07 & ~x08)))) & (~x01 | x02 | x05 | x06 | x07 | x08);
  assign n159 = ~n167 & (x07 | (n160 & ~n168 & ~n170 & n172));
  assign n160 = ~n161 & ~n164 & (n162 | ~n163) & (n165 | ~n166);
  assign n161 = ~x03 & ((~x00 & x02 & ~x06 & x08) | (x00 & ~x08 & (x02 ? (~x04 & x06) : ~x06)));
  assign n162 = (~x00 | x01 | (x02 ? (~x04 | x08) : ~x08)) & (x00 | ~x01 | x02 | ~x08);
  assign n163 = ~x03 & x06;
  assign n164 = x03 & ((~x00 & x02 & ~x04 & ~x06 & x08) | (x00 & ~x02 & x04 & x06 & ~x08));
  assign n165 = (~x00 | x01 | x06 | x08) & (x00 | ~x01 | ~x06 | ~x08);
  assign n166 = x03 & (x02 ^ ~x04);
  assign n167 = ~x03 & (x02 ? (~x06 & x07) : (x06 & (x07 | (~x00 & ~x01))));
  assign n168 = ~n169 & (x01 ? (x06 & ~x10) : (~x06 & x10));
  assign n169 = x00 ? (~x08 | (x02 ? (x03 | x04) : (~x03 | ~x04))) : (~x02 | x08 | (x03 & x04));
  assign n170 = n171 & ((~x01 & x02 & ~x05 & ~x06 & x10) | (x01 & ~x02 & x05 & x06 & ~x10));
  assign n171 = x03 & (x00 ? (~x04 & x08) : (x04 & ~x08));
  assign n172 = ~x00 | ~n126 | (x01 ? ~n174 : (~n39 | ~n173));
  assign n173 = x08 & x10;
  assign n174 = ~x10 & x08 & x06 & x04 & ~x05;
  assign n175 = x03 & ~n176;
  assign n176 = (~x07 | ((~x04 | ((x00 | ~x01 | ~x02 | ~x06) & (~x00 | ((x01 | ~x02 | ~x06) & (x02 | x06))))) & (x00 | x04 | (~x02 ^ x06)))) & (x00 | x01 | x02 | x04 | ~x06);
  assign n177 = ~n178 & n186 & (n181 | (~n182 & ~n183 & n184));
  assign n178 = ~n57 & (~n180 | (x03 & ~n179));
  assign n179 = (x01 | ~x05 | x09 | (x02 ? (x06 | ~x10) : (~x06 | x10))) & (~x01 | x02 | x05 | ~x06 | ~x09 | x10);
  assign n180 = (~x01 | x02 | ((x05 | x06 | x09) & (x03 | (~x06 ^ ~x09)))) & (x01 | ~x02 | ~x03 | ~x05 | ~x06 | ~x09);
  assign n181 = ~x06 ^ x09;
  assign n182 = ~n169 & (~x01 ^ x10);
  assign n183 = n171 & ((x05 & x10 & x01 & ~x02) | (~x01 & x02 & ~x05 & ~x10));
  assign n184 = ~x08 | (x10 ? (~n185 | ~n59) : (~n62 | ~n53));
  assign n185 = x04 & ~x05;
  assign n186 = (n189 | ~n190) & (~n59 | ~n87) & (n187 | n188);
  assign n187 = x06 ^ x09;
  assign n188 = (~x00 | ~x04 | ~x08 | (x01 ? (x02 | x03) : (~x02 | ~x03))) & (x00 | ~x01 | x02 | x04 | x08);
  assign n189 = (~x05 | ~x08 | ~x00 | x03) & (x00 | ~x03 | x05 | x08);
  assign n190 = x10 & x09 & ~x06 & x04 & x01 & x02;
  assign z07 = ~n193 | ~n209 | n216 | n222 | (~n192 & ~n206);
  assign n192 = x01 ^ x09;
  assign n193 = ~n196 & n198 & n200 & n203 & (n194 | n195);
  assign n194 = x02 ? (x03 | x04) : (~x03 | ~x04);
  assign n195 = x07 ? ((x00 | ~x08) & ((x00 & ~x08) | ((~x09 | ~x10) & (x01 | (~x09 & ~x10))))) : ((x08 | (~x00 & (~x01 | x09))) & (~x00 | ((x09 | x10) & (~x01 | (x09 & x10)))));
  assign n196 = n121 & n197 & ((x03 & ~x04 & ~x07 & ~x10) | (~x03 & x04 & (~x07 ^ x10)));
  assign n197 = x02 & ~x09;
  assign n198 = ~n199 & (~n62 | ~n30 | ~x01 | ~x02);
  assign n199 = (~x02 ^ x03) & ((~x00 & x07 & x08) | (x00 & ~x01 & ~x07 & ~x08));
  assign n200 = x00 ? (x07 | (x01 ? ~n202 : (x08 | n201))) : (~x07 | ((~x08 | n201) & (x01 | ~n202)));
  assign n201 = x02 ? (x03 | ~x04) : (~x03 | x04);
  assign n202 = ~x02 & x03 & ~x04 & ~x08;
  assign n203 = ~n204 & ((~x00 & x08) | n205 | (x00 & ~x08));
  assign n204 = ~x02 & ~x03 & ((x00 & (x01 ? (~x07 & ~x08) : (x07 & x08))) | (~x00 & ~x01 & x07 & ~x08));
  assign n205 = (~x07 | ~x09 | (x01 ? (x02 | x03) : (~x02 | (~x03 & ~x04)))) & (~x01 | x02 | x07 | x09 | (x03 & x04));
  assign n206 = (x00 | ~x02 | x08 | n207) & (~x00 | ~n69 | ~n208);
  assign n207 = x07 ? (~x10 | (~x03 ^ x04)) : x10;
  assign n208 = x10 & ~x04 & x07 & x08;
  assign n209 = (~x03 | n212) & (n210 | (~n211 & ~n215));
  assign n210 = (~x08 | (x07 ? (~x09 | ~x10) : x09)) & (x07 | ~x09 | (x08 & x10));
  assign n211 = n59 & ~x06 & x04 & x05;
  assign n212 = (x00 | ~x01 | ((x08 | n213) & (~x02 | ~n214))) & (~x00 | x01 | ~x08 | n213);
  assign n213 = (~x02 | ~x04 | x07 | x09) & (~x07 | ~x09 | x02 | x04);
  assign n214 = ~x09 & ~x08 & ~x04 & ~x07;
  assign n215 = ~x05 & x04 & ~x03 & x02 & x00 & x01;
  assign n216 = x03 & (n220 | ((x02 | ~x10) & (n217 | n218) & (~x02 | x10)));
  assign n217 = ~x08 & n51 & ((x01 & x05 & ~x07 & x09) | (~x01 & ~x05 & x07 & ~x09));
  assign n218 = n219 & ~x09 & x08 & x07 & ~x04 & ~x05;
  assign n219 = x00 & ~x01;
  assign n220 = n221 & ~x10 & x09 & x08 & x05 & ~x07;
  assign n221 = ~x04 & ~x02 & x00 & x01;
  assign n222 = x03 & (n223 | (x08 & x09 & ~x10 & n225));
  assign n223 = ~n224 & ((~x02 & ~x06 & x07 & ~x10) | (x02 & x06 & ~x07 & x10));
  assign n224 = (x00 | ~x04 | x08 | (x01 ? (x05 | ~x09) : (~x05 | x09))) & (~x00 | x01 | x04 | ~x05 | ~x08 | x09);
  assign n225 = n227 & n226 & x07 & ~x02 & ~x06;
  assign n226 = x00 & x01;
  assign n227 = ~x04 & ~x05;
  assign z08 = ~n253 | n252 | n229 | ~n236 | n242 | ~n248;
  assign n229 = x05 & (n234 | (x04 & (n230 | n233)));
  assign n230 = ~x09 & ((n146 & n232) | (x02 & ~n231));
  assign n231 = (~x00 | ~x01 | x03 | x06 | ~x08) & (~x06 | x08 | ~x10 | x00 | x01 | ~x03);
  assign n232 = ~x10 & x08 & x03 & ~x06;
  assign n233 = ~x06 & x09 & n126 & n226 & (~x08 ^ ~x10);
  assign n234 = ~n235 & n219 & ~x09 & x03 & ~x04;
  assign n235 = (~x08 | ~x10 | ~x02 | ~x06) & (x02 | x06 | x08 | x10);
  assign n236 = (n192 | n241) & (~x03 | (n237 & (~x08 | n240)));
  assign n237 = (~n221 | ~n239) & (n238 | (x02 ^ x10));
  assign n238 = (~x00 | x01 | x04 | x05 | x08 | x09) & (x00 | ~x04 | ((x08 | ~x09 | ~x01 | ~x05) & (~x08 | x09 | x01 | x05)));
  assign n239 = ~x10 & x09 & x05 & x08;
  assign n240 = (x00 | ~x01 | x02 | x04 | ~x09) & (x09 | ((x00 | x01 | x02 | x04) & (~x00 | (x01 ? (x02 | x04) : (~x02 | ~x04)))));
  assign n241 = (~x10 | ((x00 | ~x02 | ~x08 | (x03 ^ ~x04)) & (~x00 | x02 | ~x03 | x04 | x08))) & (x00 | ~x02 | x08 | x10);
  assign n242 = x03 & (n247 | (~n243 & (n244 | n246)));
  assign n243 = x02 ? (x06 | ~x10) : (~x06 | x10);
  assign n244 = ~x01 & x05 & ~x09 & ~n245;
  assign n245 = (~x00 | x04 | (x07 ^ x08)) & (x00 | ~x04 | ~x07 | x08);
  assign n246 = n40 & x07 & ~x05 & ~x00 & x01 & x04;
  assign n247 = x09 & ~x10 & n135 & n221 & (~x07 ^ x08);
  assign n248 = (n249 | ~n250) & (n251 | ((~x02 | ~x03) & n201 & (x02 | x03)));
  assign n249 = (~x00 | x02 | x04 | x06 | x08 | x10) & (x00 | ~x04 | ((x08 | ~x10 | ~x02 | ~x06) & (~x08 | x10 | x02 | x06)));
  assign n250 = x09 & ~x05 & x01 & x03;
  assign n251 = (x00 | (x01 ? (x08 | x09) : (~x08 | ~x09))) & (~x00 | x01 | x08 | ~x09);
  assign n252 = ~n194 & (x00 ? (x08 ? ((~x09 & ~x10) | (x01 & (~x09 | ~x10))) : ((x09 & x10) | (~x01 & (x09 | x10)))) : ((x01 & ~x08 & ~x09) | (x08 & ((x09 & x10) | (~x01 & (x09 | x10))))));
  assign n253 = ~n254 & ~n255 & ((~x08 & (~x09 | ~x10)) | ~n215 | (x08 & x09 & x10));
  assign n254 = ~x02 & ~x03 & (((x00 ^ x08) & (~x01 ^ x09)) | (x00 & x01 & x08 & ~x09));
  assign n255 = n219 & n197 & ((x03 & ~x04 & x08 & ~x10) | (~x03 & x04 & (~x08 ^ ~x10)));
  assign z09 = ~n272 | n281 | n283 | n285 | (~x01 & ~n257);
  assign n257 = ~n262 & ~n266 & ~n268 & (~x02 | (~n258 & n259));
  assign n258 = ~x04 & ((~x09 & ~x10 & ~x00 & x05) | (~x05 & ((~x03 & ~x09 & ~x10) | (x00 & ((~x09 & ~x10) | (x03 & x09 & x10))))));
  assign n259 = (x03 | ~x04 | ~n260) & ((~n260 & ~n261) | (x00 ? (x03 | ~x05) : (~x03 | x05)));
  assign n260 = ~x09 & ~x10;
  assign n261 = x10 & x09 & x04 & x06;
  assign n262 = n55 & ((~n263 & n265) | (x09 & ~n243 & ~n264));
  assign n263 = x02 ? (x06 | x08) : (~x06 | ~x08);
  assign n264 = (~x00 | x04 | ~x05 | x08) & (x00 | ~x04 | x05 | ~x08);
  assign n265 = ~x10 & ~x09 & ~x00 & x04 & x05;
  assign n266 = ~x10 & n69 & ~n267;
  assign n267 = (~x00 | ((x04 | ~x05 | x06 | ~x09) & (~x04 | x09))) & (x00 | ~x04 | ~x05 | x06 | ~x09);
  assign n268 = x03 & ((~n269 & n271) | (x02 & ~x06 & ~n270));
  assign n269 = ~x05 ^ x09;
  assign n270 = (~x00 | x04 | ~x05 | x07 | x09 | x10) & (x00 | ~x04 | x05 | ~x07 | ~x09 | ~x10);
  assign n271 = ~x02 & x06 & x07 & ~x10 & (x00 ^ x04);
  assign n272 = ~n277 & ~n278 & n279 & (n273 | (n70 & n274));
  assign n273 = x01 ? (~x09 ^ x10) : (~x09 | ~x10);
  assign n274 = n275 & (n263 | ~n276) & (~n135 | ~n46 | ~n69);
  assign n275 = (x00 | x02 | ~x03 | ~x04 | ~x05) & (~x00 | ((x02 | ~x03 | x04 | ~x05) & (~x02 | x03 | ~x04 | (x05 & x06))));
  assign n276 = ~x07 & ~x05 & ~x00 & x03 & x04;
  assign n277 = n72 & n28 & x10 & ~x09 & x05 & ~x08;
  assign n278 = ~x02 & (~x01 ^ ~x09) & (~x03 | (~x00 & ~x04));
  assign n279 = ~x03 | ~x04 | ((~x05 | ~x09 | ~n280) & (x09 | ~n53));
  assign n280 = ~x00 & x01 & x02;
  assign n281 = ~n282 & ~x07 & ~x00 & x03 & x04;
  assign n282 = (x05 | ((~x01 | ((~x08 | ~x09 | ~x02 | x06) & (x08 | x09 | x02 | ~x06))) & (x01 | x02 | ~x06 | x08 | ~x09))) & (x01 | ~x02 | ~x05 | x06 | ~x08 | x09);
  assign n283 = x03 & (n284 | (n185 & n280 & x06 & x09));
  assign n284 = ~n66 & ((x01 & ~x02 & ~x05 & ~x06 & ~x09) | (~x01 & ((~x06 & x09 & ~x02 & ~x05) | (x06 & ~x09 & x02 & x05))));
  assign n285 = x03 & (n287 | (x07 & ~n286 & x02 & ~x06));
  assign n286 = (x00 | ~x04 | (x01 ? (x05 | ~x09) : (~x05 | x09))) & (~x00 | x01 | x04 | ~x05 | x09);
  assign n287 = x00 & ~x02 & n72 & n227 & (~x01 ^ ~x09);
  assign z10 = n289 | ~n290 | ~n292 | ~n300 | (~x07 & ~n298);
  assign n289 = x01 & (x02 ? (~x10 & ((~x03 & ~x04) | (~x00 & (~x03 | ~x04)))) : ((x10 & (~x03 | (~x00 & ~x04))) | (x04 & ~x10 & x00 & x03)));
  assign n290 = ~n291 & (~x04 | ~x05 | x06 | x10 | ~n59);
  assign n291 = n62 & ~x10 & ~x05 & x02 & x00 & x01;
  assign n292 = ~x03 | ((~x07 | n293) & n296 & (~x10 | n297));
  assign n293 = (~x02 | x06 | ~x10 | n294) & (~x06 | x10 | ((~n227 | ~n295) & (x02 | n294)));
  assign n294 = (~x00 | x01 | x04 | ~x05) & (x00 | ~x04 | (x01 ^ ~x05));
  assign n295 = ~x02 & x00 & x01;
  assign n296 = (x00 | ~x01 | ~x02 | ~x04 | ~x05 | ~x10) & ((~x00 ^ x04) | ((x01 | x05 | (~x02 ^ x10)) & (~x01 | x02 | ~x05 | x10)));
  assign n297 = (~x04 & (~x00 | (~x05 & x06))) | (~x02 & x06) | (~x01 & ~x05) | (x00 & x04) | (x02 & ~x06) | (x01 & x05);
  assign n298 = (~n171 | n299) & (x08 | ~n28 | ~n29 | ~n260);
  assign n299 = (~x01 | x02 | x05 | ~x06 | x09 | ~x10) & (x01 | ~x05 | ((~x02 | x06 | (~x09 ^ ~x10)) & (~x09 | x10 | x02 | ~x06)));
  assign n300 = (x01 | (n301 & (~x05 | ~n55 | n302))) & (~x01 | x05 | ~n55 | n303);
  assign n301 = (~x00 | ~x03 | ~x04 | (~x02 ^ ~x10)) & ((x02 ^ ~x10) | (x03 & (x00 | x04)));
  assign n302 = x00 ? (x04 | x08 | (x02 ? (x06 | x10) : (~x06 | ~x10))) : (~x04 | ~x08 | (x02 ? (x06 | ~x10) : (~x06 | x10)));
  assign n303 = (~x00 | x02 | x04 | ~x06 | x08 | ~x10) & (x00 | ~x04 | ((~x02 | x06 | (~x08 ^ ~x10)) & (~x08 | x10 | x02 | ~x06)));
endmodule


