module div_24_241(X, Q, R );

input  [24:1] X;
output [17:1] Q;  
output [8:1] R;  

wire [17:1] Q_temp;
wire [10:1] r_1;
wire [9:1] r_2;
wire r_3;

wire [10:1] sum_res;
wire [10:1] sum;

wire [17:1] q_1;
wire [25:1] q_2;

q_1 label1 ( .x0(X[16]),.x1(X[15]),.x2(X[14]),.x3(X[13]),.x4(X[12]),.x5(X[11]),.x6(X[10]),.x7(X[9]),
.z00(q_1[17]),.z01(q_1[16]),.z02(q_1[15]),.z03(q_1[14]),.z04(q_1[13]),.z05(q_1[12]),.z06(q_1[11]),.z07(q_1[10]),.z08(q_1[9]),.z09(q_1[8]),.z10(q_1[7]),.z11(q_1[6]),.z12(q_1[5]),.z13(q_1[4]),.z14(q_1[3]),.z15(q_1[2]),.z16(q_1[1]));

q_2 label2 ( .x0(X[24]),.x1(X[23]),.x2(X[22]),.x3(X[21]),.x4(X[20]),.x5(X[19]),.x6(X[18]),.x7(X[17]),
.z00(q_2[25]),.z01(q_2[24]),.z02(q_2[23]),.z03(q_2[22]),.z04(q_2[21]),.z05(q_2[20]),.z06(q_2[19]),.z07(q_2[18]),.z08(q_2[17]),.z09(q_2[16]),.z10(q_2[15]),.z11(q_2[14]),.z12(q_2[13]),.z13(q_2[12]),.z14(q_2[11]),.z15(q_2[10]),.z16(q_2[9]),.z17(q_2[8]),.z18(q_2[7]),.z19(q_2[6]),.z20(q_2[5]),.z21(q_2[4]),.z22(q_2[3]),.z23(q_2[2]),.z24(q_2[1]));


assign sum_res = X[8:1] + q_1[8:1] + q_2[8:1];

quot_res  label8 (.x0(sum_res[10]),.x1(sum_res[9]),.x2(sum_res[8]),.x3(sum_res[7]),.x4(sum_res[6]),.x5(sum_res[5]),.x6(sum_res[4]),
		  .x7(sum_res[3]),.x8(sum_res[2]),.x9(sum_res[1]),
                  .z0(sum[10]),.z1(sum[9]),.z2(sum[8]),.z3(sum[7]),.z4(sum[6]),.z5(sum[5]),.z6(sum[4]),
		  .z7(sum[3]),.z8(sum[2]),.z9(sum[1]));

assign r_1 = q_1[16:9] + q_2[16:9];

assign r_2 = q_1[17] + r_1[9] + q_2[24:17];

assign r_3 = q_2[25];

assign Q_temp = {r_3, r_2[8:1], r_1[8:1]};


assign Q = Q_temp + sum[10:9];

assign R = sum[8:1]; 

endmodule