// Benchmark "q_3" written by ABC on Mon Jul 10 22:15:59 2023

module q_3 ( 
    x0,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15  );
  input  x0;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15;
  assign z00 = x0;
  assign z01 = x0;
  assign z02 = 1'b0;
  assign z03 = 1'b0;
  assign z04 = x0;
  assign z05 = x0;
  assign z06 = 1'b0;
  assign z07 = 1'b0;
  assign z08 = x0;
  assign z09 = x0;
  assign z10 = 1'b0;
  assign z11 = 1'b0;
  assign z12 = x0;
  assign z13 = 1'b0;
  assign z14 = x0;
  assign z15 = x0;
endmodule


