module div_24_113(X, Q, R );

input  [24:1] X;
output [18:1] Q;  
output [7:1] R;  

wire [18:1] Q_temp;
wire [9:1] r_1;
wire [8:1] r_2;
wire [4:1] r_3;

wire [9:1] sum_res;
wire [10:1] sum;

wire [15:1] q_1;
wire [22:1] q_2;
wire [25:1] q_3;

q_1 label1 ( .x0(X[14]),.x1(X[13]),.x2(X[12]),.x3(X[11]),.x4(X[10]),.x5(X[9]),.x6(X[8]),
.z00(q_1[15]),.z01(q_1[14]),.z02(q_1[13]),.z03(q_1[12]),.z04(q_1[11]),.z05(q_1[10]),.z06(q_1[9]),.z07(q_1[8]),.z08(q_1[7]),.z09(q_1[6]),.z10(q_1[5]),.z11(q_1[4]),.z12(q_1[3]),.z13(q_1[2]),.z14(q_1[1]));

q_2 label2 ( .x0(X[21]),.x1(X[20]),.x2(X[19]),.x3(X[18]),.x4(X[17]),.x5(X[16]),.x6(X[15]),
.z00(q_2[22]),.z01(q_2[21]),.z02(q_2[20]),.z03(q_2[19]),.z04(q_2[18]),.z05(q_2[17]),.z06(q_2[16]),.z07(q_2[15]),.z08(q_2[14]),.z09(q_2[13]),.z10(q_2[12]),.z11(q_2[11]),.z12(q_2[10]),.z13(q_2[9]),.z14(q_2[8]),.z15(q_2[7]),.z16(q_2[6]),.z17(q_2[5]),.z18(q_2[4]),.z19(q_2[3]),.z20(q_2[2]),.z21(q_2[1]));

q_3 label3 ( .x0(X[24]),.x1(X[23]),.x2(X[22]),
.z00(q_3[24]),.z01(q_3[23]),.z02(q_3[22]),.z03(q_3[21]),.z04(q_3[20]),.z05(q_3[19]),.z06(q_3[18]),.z07(q_3[17]),.z08(q_3[16]),.z09(q_3[15]),.z10(q_3[14]),.z11(q_3[13]),.z12(q_3[12]),.z13(q_3[11]),.z14(q_3[10]),.z15(q_3[9]),.z16(q_3[8]),.z17(q_3[7]),.z18(q_3[6]),.z19(q_3[5]),.z20(q_3[4]),.z21(q_3[3]),.z22(q_3[2]),.z23(q_3[1]));


assign sum_res = X[7:1] + q_1[7:1] + q_2[7:1] + q_3[7:1];

quot_res  label9 (.x0(sum_res[9]),.x1(sum_res[8]),.x2(sum_res[7]),.x3(sum_res[6]),.x4(sum_res[5]),.x5(sum_res[4]),
		  .x6(sum_res[3]),.x7(sum_res[2]),.x8(sum_res[1]),
                  .z0(sum[10]),.z1(sum[9]),.z2(sum[8]),.z3(sum[7]),.z4(sum[6]),.z5(sum[5]),
		  .z6(sum[4]),.z7(sum[3]),.z8(sum[2]),.z9(sum[1]));

assign r_1 = q_1[14:8] + q_2[14:8] + q_3[14:8];

assign r_2 = q_1[15] + r_1[9:8] + q_2[21:15] + q_3[21:15];

assign r_3 = r_2[8] + q_2[22] + q_3[24:22];


assign Q_temp = {r_3[4:1], r_2[7:1], r_1[7:1]};

assign Q = Q_temp + sum[10:8];

assign R = sum[7:1]; 

endmodule