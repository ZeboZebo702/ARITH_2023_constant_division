// Benchmark "q_3" written by ABC on Mon Jul 10 22:36:39 2023

module q_3 ( 
    x0,
    z0, z1, z2  );
  input  x0;
  output z0, z1, z2;
  assign z0 = 1'b0;
  assign z1 = x0;
  assign z2 = x0;
endmodule


