// Benchmark "q_11" written by ABC on Tue Jul 11 01:37:07 2023

module q_11 ( 
    x0,
    z0, z1, z2  );
  input  x0;
  output z0, z1, z2;
  assign z0 = 1'b0;
  assign z1 = x0;
  assign z2 = x0;
endmodule


